magic
tech gf180mcuD
magscale 1 5
timestamp 1701352414
<< obsm1 >>
rect 672 1471 299320 298577
<< metal2 >>
rect 2128 299600 2184 300000
rect 4368 299600 4424 300000
rect 6608 299600 6664 300000
rect 8848 299600 8904 300000
rect 11088 299600 11144 300000
rect 13328 299600 13384 300000
rect 15568 299600 15624 300000
rect 17808 299600 17864 300000
rect 20048 299600 20104 300000
rect 22288 299600 22344 300000
rect 24528 299600 24584 300000
rect 26768 299600 26824 300000
rect 29008 299600 29064 300000
rect 31248 299600 31304 300000
rect 33488 299600 33544 300000
rect 35728 299600 35784 300000
rect 37968 299600 38024 300000
rect 40208 299600 40264 300000
rect 42448 299600 42504 300000
rect 44688 299600 44744 300000
rect 46928 299600 46984 300000
rect 49168 299600 49224 300000
rect 51408 299600 51464 300000
rect 53648 299600 53704 300000
rect 55888 299600 55944 300000
rect 58128 299600 58184 300000
rect 60368 299600 60424 300000
rect 62608 299600 62664 300000
rect 64848 299600 64904 300000
rect 67088 299600 67144 300000
rect 69328 299600 69384 300000
rect 71568 299600 71624 300000
rect 73808 299600 73864 300000
rect 76048 299600 76104 300000
rect 78288 299600 78344 300000
rect 80528 299600 80584 300000
rect 82768 299600 82824 300000
rect 85008 299600 85064 300000
rect 87248 299600 87304 300000
rect 89488 299600 89544 300000
rect 91728 299600 91784 300000
rect 93968 299600 94024 300000
rect 96208 299600 96264 300000
rect 98448 299600 98504 300000
rect 100688 299600 100744 300000
rect 102928 299600 102984 300000
rect 105168 299600 105224 300000
rect 107408 299600 107464 300000
rect 109648 299600 109704 300000
rect 111888 299600 111944 300000
rect 114128 299600 114184 300000
rect 116368 299600 116424 300000
rect 118608 299600 118664 300000
rect 120848 299600 120904 300000
rect 123088 299600 123144 300000
rect 125328 299600 125384 300000
rect 127568 299600 127624 300000
rect 129808 299600 129864 300000
rect 132048 299600 132104 300000
rect 134288 299600 134344 300000
rect 136528 299600 136584 300000
rect 138768 299600 138824 300000
rect 141008 299600 141064 300000
rect 143248 299600 143304 300000
rect 145488 299600 145544 300000
rect 147728 299600 147784 300000
rect 149968 299600 150024 300000
rect 152208 299600 152264 300000
rect 154448 299600 154504 300000
rect 156688 299600 156744 300000
rect 158928 299600 158984 300000
rect 161168 299600 161224 300000
rect 163408 299600 163464 300000
rect 165648 299600 165704 300000
rect 167888 299600 167944 300000
rect 170128 299600 170184 300000
rect 172368 299600 172424 300000
rect 174608 299600 174664 300000
rect 176848 299600 176904 300000
rect 179088 299600 179144 300000
rect 181328 299600 181384 300000
rect 183568 299600 183624 300000
rect 185808 299600 185864 300000
rect 188048 299600 188104 300000
rect 190288 299600 190344 300000
rect 192528 299600 192584 300000
rect 194768 299600 194824 300000
rect 197008 299600 197064 300000
rect 199248 299600 199304 300000
rect 201488 299600 201544 300000
rect 203728 299600 203784 300000
rect 205968 299600 206024 300000
rect 208208 299600 208264 300000
rect 210448 299600 210504 300000
rect 212688 299600 212744 300000
rect 214928 299600 214984 300000
rect 217168 299600 217224 300000
rect 219408 299600 219464 300000
rect 221648 299600 221704 300000
rect 223888 299600 223944 300000
rect 226128 299600 226184 300000
rect 228368 299600 228424 300000
rect 230608 299600 230664 300000
rect 232848 299600 232904 300000
rect 235088 299600 235144 300000
rect 237328 299600 237384 300000
rect 239568 299600 239624 300000
rect 241808 299600 241864 300000
rect 244048 299600 244104 300000
rect 246288 299600 246344 300000
rect 248528 299600 248584 300000
rect 250768 299600 250824 300000
rect 253008 299600 253064 300000
rect 255248 299600 255304 300000
rect 257488 299600 257544 300000
rect 259728 299600 259784 300000
rect 261968 299600 262024 300000
rect 264208 299600 264264 300000
rect 266448 299600 266504 300000
rect 268688 299600 268744 300000
rect 270928 299600 270984 300000
rect 273168 299600 273224 300000
rect 275408 299600 275464 300000
rect 277648 299600 277704 300000
rect 279888 299600 279944 300000
rect 282128 299600 282184 300000
rect 284368 299600 284424 300000
rect 286608 299600 286664 300000
rect 288848 299600 288904 300000
rect 291088 299600 291144 300000
rect 293328 299600 293384 300000
rect 295568 299600 295624 300000
rect 297808 299600 297864 300000
rect 13328 0 13384 400
rect 14448 0 14504 400
rect 15568 0 15624 400
rect 16688 0 16744 400
rect 17808 0 17864 400
rect 18928 0 18984 400
rect 20048 0 20104 400
rect 21168 0 21224 400
rect 22288 0 22344 400
rect 23408 0 23464 400
rect 24528 0 24584 400
rect 25648 0 25704 400
rect 26768 0 26824 400
rect 27888 0 27944 400
rect 29008 0 29064 400
rect 30128 0 30184 400
rect 31248 0 31304 400
rect 32368 0 32424 400
rect 33488 0 33544 400
rect 34608 0 34664 400
rect 35728 0 35784 400
rect 36848 0 36904 400
rect 37968 0 38024 400
rect 39088 0 39144 400
rect 40208 0 40264 400
rect 41328 0 41384 400
rect 42448 0 42504 400
rect 43568 0 43624 400
rect 44688 0 44744 400
rect 45808 0 45864 400
rect 46928 0 46984 400
rect 48048 0 48104 400
rect 49168 0 49224 400
rect 50288 0 50344 400
rect 51408 0 51464 400
rect 52528 0 52584 400
rect 53648 0 53704 400
rect 54768 0 54824 400
rect 55888 0 55944 400
rect 57008 0 57064 400
rect 58128 0 58184 400
rect 59248 0 59304 400
rect 60368 0 60424 400
rect 61488 0 61544 400
rect 62608 0 62664 400
rect 63728 0 63784 400
rect 64848 0 64904 400
rect 65968 0 66024 400
rect 67088 0 67144 400
rect 68208 0 68264 400
rect 69328 0 69384 400
rect 70448 0 70504 400
rect 71568 0 71624 400
rect 72688 0 72744 400
rect 73808 0 73864 400
rect 74928 0 74984 400
rect 76048 0 76104 400
rect 77168 0 77224 400
rect 78288 0 78344 400
rect 79408 0 79464 400
rect 80528 0 80584 400
rect 81648 0 81704 400
rect 82768 0 82824 400
rect 83888 0 83944 400
rect 85008 0 85064 400
rect 86128 0 86184 400
rect 87248 0 87304 400
rect 88368 0 88424 400
rect 89488 0 89544 400
rect 90608 0 90664 400
rect 91728 0 91784 400
rect 92848 0 92904 400
rect 93968 0 94024 400
rect 95088 0 95144 400
rect 96208 0 96264 400
rect 97328 0 97384 400
rect 98448 0 98504 400
rect 99568 0 99624 400
rect 100688 0 100744 400
rect 101808 0 101864 400
rect 102928 0 102984 400
rect 104048 0 104104 400
rect 105168 0 105224 400
rect 106288 0 106344 400
rect 107408 0 107464 400
rect 108528 0 108584 400
rect 109648 0 109704 400
rect 110768 0 110824 400
rect 111888 0 111944 400
rect 113008 0 113064 400
rect 114128 0 114184 400
rect 115248 0 115304 400
rect 116368 0 116424 400
rect 117488 0 117544 400
rect 118608 0 118664 400
rect 119728 0 119784 400
rect 120848 0 120904 400
rect 121968 0 122024 400
rect 123088 0 123144 400
rect 124208 0 124264 400
rect 125328 0 125384 400
rect 126448 0 126504 400
rect 127568 0 127624 400
rect 128688 0 128744 400
rect 129808 0 129864 400
rect 130928 0 130984 400
rect 132048 0 132104 400
rect 133168 0 133224 400
rect 134288 0 134344 400
rect 135408 0 135464 400
rect 136528 0 136584 400
rect 137648 0 137704 400
rect 138768 0 138824 400
rect 139888 0 139944 400
rect 141008 0 141064 400
rect 142128 0 142184 400
rect 143248 0 143304 400
rect 144368 0 144424 400
rect 145488 0 145544 400
rect 146608 0 146664 400
rect 147728 0 147784 400
rect 148848 0 148904 400
rect 149968 0 150024 400
rect 151088 0 151144 400
rect 152208 0 152264 400
rect 153328 0 153384 400
rect 154448 0 154504 400
rect 155568 0 155624 400
rect 156688 0 156744 400
rect 157808 0 157864 400
rect 158928 0 158984 400
rect 160048 0 160104 400
rect 161168 0 161224 400
rect 162288 0 162344 400
rect 163408 0 163464 400
rect 164528 0 164584 400
rect 165648 0 165704 400
rect 166768 0 166824 400
rect 167888 0 167944 400
rect 169008 0 169064 400
rect 170128 0 170184 400
rect 171248 0 171304 400
rect 172368 0 172424 400
rect 173488 0 173544 400
rect 174608 0 174664 400
rect 175728 0 175784 400
rect 176848 0 176904 400
rect 177968 0 178024 400
rect 179088 0 179144 400
rect 180208 0 180264 400
rect 181328 0 181384 400
rect 182448 0 182504 400
rect 183568 0 183624 400
rect 184688 0 184744 400
rect 185808 0 185864 400
rect 186928 0 186984 400
rect 188048 0 188104 400
rect 189168 0 189224 400
rect 190288 0 190344 400
rect 191408 0 191464 400
rect 192528 0 192584 400
rect 193648 0 193704 400
rect 194768 0 194824 400
rect 195888 0 195944 400
rect 197008 0 197064 400
rect 198128 0 198184 400
rect 199248 0 199304 400
rect 200368 0 200424 400
rect 201488 0 201544 400
rect 202608 0 202664 400
rect 203728 0 203784 400
rect 204848 0 204904 400
rect 205968 0 206024 400
rect 207088 0 207144 400
rect 208208 0 208264 400
rect 209328 0 209384 400
rect 210448 0 210504 400
rect 211568 0 211624 400
rect 212688 0 212744 400
rect 213808 0 213864 400
rect 214928 0 214984 400
rect 216048 0 216104 400
rect 217168 0 217224 400
rect 218288 0 218344 400
rect 219408 0 219464 400
rect 220528 0 220584 400
rect 221648 0 221704 400
rect 222768 0 222824 400
rect 223888 0 223944 400
rect 225008 0 225064 400
rect 226128 0 226184 400
rect 227248 0 227304 400
rect 228368 0 228424 400
rect 229488 0 229544 400
rect 230608 0 230664 400
rect 231728 0 231784 400
rect 232848 0 232904 400
rect 233968 0 234024 400
rect 235088 0 235144 400
rect 236208 0 236264 400
rect 237328 0 237384 400
rect 238448 0 238504 400
rect 239568 0 239624 400
rect 240688 0 240744 400
rect 241808 0 241864 400
rect 242928 0 242984 400
rect 244048 0 244104 400
rect 245168 0 245224 400
rect 246288 0 246344 400
rect 247408 0 247464 400
rect 248528 0 248584 400
rect 249648 0 249704 400
rect 250768 0 250824 400
rect 251888 0 251944 400
rect 253008 0 253064 400
rect 254128 0 254184 400
rect 255248 0 255304 400
rect 256368 0 256424 400
rect 257488 0 257544 400
rect 258608 0 258664 400
rect 259728 0 259784 400
rect 260848 0 260904 400
rect 261968 0 262024 400
rect 263088 0 263144 400
rect 264208 0 264264 400
rect 265328 0 265384 400
rect 266448 0 266504 400
rect 267568 0 267624 400
rect 268688 0 268744 400
rect 269808 0 269864 400
rect 270928 0 270984 400
rect 272048 0 272104 400
rect 273168 0 273224 400
rect 274288 0 274344 400
rect 275408 0 275464 400
rect 276528 0 276584 400
rect 277648 0 277704 400
rect 278768 0 278824 400
rect 279888 0 279944 400
rect 281008 0 281064 400
rect 282128 0 282184 400
rect 283248 0 283304 400
rect 284368 0 284424 400
rect 285488 0 285544 400
rect 286608 0 286664 400
<< obsm2 >>
rect 14 299570 2098 299983
rect 2214 299570 4338 299983
rect 4454 299570 6578 299983
rect 6694 299570 8818 299983
rect 8934 299570 11058 299983
rect 11174 299570 13298 299983
rect 13414 299570 15538 299983
rect 15654 299570 17778 299983
rect 17894 299570 20018 299983
rect 20134 299570 22258 299983
rect 22374 299570 24498 299983
rect 24614 299570 26738 299983
rect 26854 299570 28978 299983
rect 29094 299570 31218 299983
rect 31334 299570 33458 299983
rect 33574 299570 35698 299983
rect 35814 299570 37938 299983
rect 38054 299570 40178 299983
rect 40294 299570 42418 299983
rect 42534 299570 44658 299983
rect 44774 299570 46898 299983
rect 47014 299570 49138 299983
rect 49254 299570 51378 299983
rect 51494 299570 53618 299983
rect 53734 299570 55858 299983
rect 55974 299570 58098 299983
rect 58214 299570 60338 299983
rect 60454 299570 62578 299983
rect 62694 299570 64818 299983
rect 64934 299570 67058 299983
rect 67174 299570 69298 299983
rect 69414 299570 71538 299983
rect 71654 299570 73778 299983
rect 73894 299570 76018 299983
rect 76134 299570 78258 299983
rect 78374 299570 80498 299983
rect 80614 299570 82738 299983
rect 82854 299570 84978 299983
rect 85094 299570 87218 299983
rect 87334 299570 89458 299983
rect 89574 299570 91698 299983
rect 91814 299570 93938 299983
rect 94054 299570 96178 299983
rect 96294 299570 98418 299983
rect 98534 299570 100658 299983
rect 100774 299570 102898 299983
rect 103014 299570 105138 299983
rect 105254 299570 107378 299983
rect 107494 299570 109618 299983
rect 109734 299570 111858 299983
rect 111974 299570 114098 299983
rect 114214 299570 116338 299983
rect 116454 299570 118578 299983
rect 118694 299570 120818 299983
rect 120934 299570 123058 299983
rect 123174 299570 125298 299983
rect 125414 299570 127538 299983
rect 127654 299570 129778 299983
rect 129894 299570 132018 299983
rect 132134 299570 134258 299983
rect 134374 299570 136498 299983
rect 136614 299570 138738 299983
rect 138854 299570 140978 299983
rect 141094 299570 143218 299983
rect 143334 299570 145458 299983
rect 145574 299570 147698 299983
rect 147814 299570 149938 299983
rect 150054 299570 152178 299983
rect 152294 299570 154418 299983
rect 154534 299570 156658 299983
rect 156774 299570 158898 299983
rect 159014 299570 161138 299983
rect 161254 299570 163378 299983
rect 163494 299570 165618 299983
rect 165734 299570 167858 299983
rect 167974 299570 170098 299983
rect 170214 299570 172338 299983
rect 172454 299570 174578 299983
rect 174694 299570 176818 299983
rect 176934 299570 179058 299983
rect 179174 299570 181298 299983
rect 181414 299570 183538 299983
rect 183654 299570 185778 299983
rect 185894 299570 188018 299983
rect 188134 299570 190258 299983
rect 190374 299570 192498 299983
rect 192614 299570 194738 299983
rect 194854 299570 196978 299983
rect 197094 299570 199218 299983
rect 199334 299570 201458 299983
rect 201574 299570 203698 299983
rect 203814 299570 205938 299983
rect 206054 299570 208178 299983
rect 208294 299570 210418 299983
rect 210534 299570 212658 299983
rect 212774 299570 214898 299983
rect 215014 299570 217138 299983
rect 217254 299570 219378 299983
rect 219494 299570 221618 299983
rect 221734 299570 223858 299983
rect 223974 299570 226098 299983
rect 226214 299570 228338 299983
rect 228454 299570 230578 299983
rect 230694 299570 232818 299983
rect 232934 299570 235058 299983
rect 235174 299570 237298 299983
rect 237414 299570 239538 299983
rect 239654 299570 241778 299983
rect 241894 299570 244018 299983
rect 244134 299570 246258 299983
rect 246374 299570 248498 299983
rect 248614 299570 250738 299983
rect 250854 299570 252978 299983
rect 253094 299570 255218 299983
rect 255334 299570 257458 299983
rect 257574 299570 259698 299983
rect 259814 299570 261938 299983
rect 262054 299570 264178 299983
rect 264294 299570 266418 299983
rect 266534 299570 268658 299983
rect 268774 299570 270898 299983
rect 271014 299570 273138 299983
rect 273254 299570 275378 299983
rect 275494 299570 277618 299983
rect 277734 299570 279858 299983
rect 279974 299570 282098 299983
rect 282214 299570 284338 299983
rect 284454 299570 286578 299983
rect 286694 299570 288818 299983
rect 288934 299570 291058 299983
rect 291174 299570 293298 299983
rect 293414 299570 295538 299983
rect 295654 299570 297778 299983
rect 297894 299570 299362 299983
rect 14 430 299362 299570
rect 14 9 13298 430
rect 13414 9 14418 430
rect 14534 9 15538 430
rect 15654 9 16658 430
rect 16774 9 17778 430
rect 17894 9 18898 430
rect 19014 9 20018 430
rect 20134 9 21138 430
rect 21254 9 22258 430
rect 22374 9 23378 430
rect 23494 9 24498 430
rect 24614 9 25618 430
rect 25734 9 26738 430
rect 26854 9 27858 430
rect 27974 9 28978 430
rect 29094 9 30098 430
rect 30214 9 31218 430
rect 31334 9 32338 430
rect 32454 9 33458 430
rect 33574 9 34578 430
rect 34694 9 35698 430
rect 35814 9 36818 430
rect 36934 9 37938 430
rect 38054 9 39058 430
rect 39174 9 40178 430
rect 40294 9 41298 430
rect 41414 9 42418 430
rect 42534 9 43538 430
rect 43654 9 44658 430
rect 44774 9 45778 430
rect 45894 9 46898 430
rect 47014 9 48018 430
rect 48134 9 49138 430
rect 49254 9 50258 430
rect 50374 9 51378 430
rect 51494 9 52498 430
rect 52614 9 53618 430
rect 53734 9 54738 430
rect 54854 9 55858 430
rect 55974 9 56978 430
rect 57094 9 58098 430
rect 58214 9 59218 430
rect 59334 9 60338 430
rect 60454 9 61458 430
rect 61574 9 62578 430
rect 62694 9 63698 430
rect 63814 9 64818 430
rect 64934 9 65938 430
rect 66054 9 67058 430
rect 67174 9 68178 430
rect 68294 9 69298 430
rect 69414 9 70418 430
rect 70534 9 71538 430
rect 71654 9 72658 430
rect 72774 9 73778 430
rect 73894 9 74898 430
rect 75014 9 76018 430
rect 76134 9 77138 430
rect 77254 9 78258 430
rect 78374 9 79378 430
rect 79494 9 80498 430
rect 80614 9 81618 430
rect 81734 9 82738 430
rect 82854 9 83858 430
rect 83974 9 84978 430
rect 85094 9 86098 430
rect 86214 9 87218 430
rect 87334 9 88338 430
rect 88454 9 89458 430
rect 89574 9 90578 430
rect 90694 9 91698 430
rect 91814 9 92818 430
rect 92934 9 93938 430
rect 94054 9 95058 430
rect 95174 9 96178 430
rect 96294 9 97298 430
rect 97414 9 98418 430
rect 98534 9 99538 430
rect 99654 9 100658 430
rect 100774 9 101778 430
rect 101894 9 102898 430
rect 103014 9 104018 430
rect 104134 9 105138 430
rect 105254 9 106258 430
rect 106374 9 107378 430
rect 107494 9 108498 430
rect 108614 9 109618 430
rect 109734 9 110738 430
rect 110854 9 111858 430
rect 111974 9 112978 430
rect 113094 9 114098 430
rect 114214 9 115218 430
rect 115334 9 116338 430
rect 116454 9 117458 430
rect 117574 9 118578 430
rect 118694 9 119698 430
rect 119814 9 120818 430
rect 120934 9 121938 430
rect 122054 9 123058 430
rect 123174 9 124178 430
rect 124294 9 125298 430
rect 125414 9 126418 430
rect 126534 9 127538 430
rect 127654 9 128658 430
rect 128774 9 129778 430
rect 129894 9 130898 430
rect 131014 9 132018 430
rect 132134 9 133138 430
rect 133254 9 134258 430
rect 134374 9 135378 430
rect 135494 9 136498 430
rect 136614 9 137618 430
rect 137734 9 138738 430
rect 138854 9 139858 430
rect 139974 9 140978 430
rect 141094 9 142098 430
rect 142214 9 143218 430
rect 143334 9 144338 430
rect 144454 9 145458 430
rect 145574 9 146578 430
rect 146694 9 147698 430
rect 147814 9 148818 430
rect 148934 9 149938 430
rect 150054 9 151058 430
rect 151174 9 152178 430
rect 152294 9 153298 430
rect 153414 9 154418 430
rect 154534 9 155538 430
rect 155654 9 156658 430
rect 156774 9 157778 430
rect 157894 9 158898 430
rect 159014 9 160018 430
rect 160134 9 161138 430
rect 161254 9 162258 430
rect 162374 9 163378 430
rect 163494 9 164498 430
rect 164614 9 165618 430
rect 165734 9 166738 430
rect 166854 9 167858 430
rect 167974 9 168978 430
rect 169094 9 170098 430
rect 170214 9 171218 430
rect 171334 9 172338 430
rect 172454 9 173458 430
rect 173574 9 174578 430
rect 174694 9 175698 430
rect 175814 9 176818 430
rect 176934 9 177938 430
rect 178054 9 179058 430
rect 179174 9 180178 430
rect 180294 9 181298 430
rect 181414 9 182418 430
rect 182534 9 183538 430
rect 183654 9 184658 430
rect 184774 9 185778 430
rect 185894 9 186898 430
rect 187014 9 188018 430
rect 188134 9 189138 430
rect 189254 9 190258 430
rect 190374 9 191378 430
rect 191494 9 192498 430
rect 192614 9 193618 430
rect 193734 9 194738 430
rect 194854 9 195858 430
rect 195974 9 196978 430
rect 197094 9 198098 430
rect 198214 9 199218 430
rect 199334 9 200338 430
rect 200454 9 201458 430
rect 201574 9 202578 430
rect 202694 9 203698 430
rect 203814 9 204818 430
rect 204934 9 205938 430
rect 206054 9 207058 430
rect 207174 9 208178 430
rect 208294 9 209298 430
rect 209414 9 210418 430
rect 210534 9 211538 430
rect 211654 9 212658 430
rect 212774 9 213778 430
rect 213894 9 214898 430
rect 215014 9 216018 430
rect 216134 9 217138 430
rect 217254 9 218258 430
rect 218374 9 219378 430
rect 219494 9 220498 430
rect 220614 9 221618 430
rect 221734 9 222738 430
rect 222854 9 223858 430
rect 223974 9 224978 430
rect 225094 9 226098 430
rect 226214 9 227218 430
rect 227334 9 228338 430
rect 228454 9 229458 430
rect 229574 9 230578 430
rect 230694 9 231698 430
rect 231814 9 232818 430
rect 232934 9 233938 430
rect 234054 9 235058 430
rect 235174 9 236178 430
rect 236294 9 237298 430
rect 237414 9 238418 430
rect 238534 9 239538 430
rect 239654 9 240658 430
rect 240774 9 241778 430
rect 241894 9 242898 430
rect 243014 9 244018 430
rect 244134 9 245138 430
rect 245254 9 246258 430
rect 246374 9 247378 430
rect 247494 9 248498 430
rect 248614 9 249618 430
rect 249734 9 250738 430
rect 250854 9 251858 430
rect 251974 9 252978 430
rect 253094 9 254098 430
rect 254214 9 255218 430
rect 255334 9 256338 430
rect 256454 9 257458 430
rect 257574 9 258578 430
rect 258694 9 259698 430
rect 259814 9 260818 430
rect 260934 9 261938 430
rect 262054 9 263058 430
rect 263174 9 264178 430
rect 264294 9 265298 430
rect 265414 9 266418 430
rect 266534 9 267538 430
rect 267654 9 268658 430
rect 268774 9 269778 430
rect 269894 9 270898 430
rect 271014 9 272018 430
rect 272134 9 273138 430
rect 273254 9 274258 430
rect 274374 9 275378 430
rect 275494 9 276498 430
rect 276614 9 277618 430
rect 277734 9 278738 430
rect 278854 9 279858 430
rect 279974 9 280978 430
rect 281094 9 282098 430
rect 282214 9 283218 430
rect 283334 9 284338 430
rect 284454 9 285458 430
rect 285574 9 286578 430
rect 286694 9 299362 430
<< metal3 >>
rect 0 294448 400 294504
rect 0 292208 400 292264
rect 0 289968 400 290024
rect 0 287728 400 287784
rect 0 285488 400 285544
rect 0 283248 400 283304
rect 0 281008 400 281064
rect 0 278768 400 278824
rect 0 276528 400 276584
rect 0 274288 400 274344
rect 0 272048 400 272104
rect 0 269808 400 269864
rect 0 267568 400 267624
rect 0 265328 400 265384
rect 0 263088 400 263144
rect 0 260848 400 260904
rect 0 258608 400 258664
rect 0 256368 400 256424
rect 0 254128 400 254184
rect 0 251888 400 251944
rect 0 249648 400 249704
rect 0 247408 400 247464
rect 0 245168 400 245224
rect 0 242928 400 242984
rect 0 240688 400 240744
rect 0 238448 400 238504
rect 0 236208 400 236264
rect 0 233968 400 234024
rect 0 231728 400 231784
rect 0 229488 400 229544
rect 0 227248 400 227304
rect 0 225008 400 225064
rect 0 222768 400 222824
rect 0 220528 400 220584
rect 0 218288 400 218344
rect 0 216048 400 216104
rect 0 213808 400 213864
rect 0 211568 400 211624
rect 0 209328 400 209384
rect 0 207088 400 207144
rect 0 204848 400 204904
rect 0 202608 400 202664
rect 0 200368 400 200424
rect 0 198128 400 198184
rect 0 195888 400 195944
rect 0 193648 400 193704
rect 0 191408 400 191464
rect 0 189168 400 189224
rect 0 186928 400 186984
rect 0 184688 400 184744
rect 0 182448 400 182504
rect 0 180208 400 180264
rect 0 177968 400 178024
rect 0 175728 400 175784
rect 0 173488 400 173544
rect 0 171248 400 171304
rect 0 169008 400 169064
rect 0 166768 400 166824
rect 0 164528 400 164584
rect 0 162288 400 162344
rect 0 160048 400 160104
rect 0 157808 400 157864
rect 0 155568 400 155624
rect 0 153328 400 153384
rect 0 151088 400 151144
rect 0 148848 400 148904
rect 0 146608 400 146664
rect 0 144368 400 144424
rect 0 142128 400 142184
rect 0 139888 400 139944
rect 0 137648 400 137704
rect 0 135408 400 135464
rect 0 133168 400 133224
rect 0 130928 400 130984
rect 0 128688 400 128744
rect 0 126448 400 126504
rect 0 124208 400 124264
rect 0 121968 400 122024
rect 0 119728 400 119784
rect 0 117488 400 117544
rect 0 115248 400 115304
rect 0 113008 400 113064
rect 0 110768 400 110824
rect 0 108528 400 108584
rect 0 106288 400 106344
rect 0 104048 400 104104
rect 0 101808 400 101864
rect 0 99568 400 99624
rect 0 97328 400 97384
rect 0 95088 400 95144
rect 0 92848 400 92904
rect 0 90608 400 90664
rect 0 88368 400 88424
rect 0 86128 400 86184
rect 0 83888 400 83944
rect 0 81648 400 81704
rect 0 79408 400 79464
rect 0 77168 400 77224
rect 0 74928 400 74984
rect 0 72688 400 72744
rect 0 70448 400 70504
rect 0 68208 400 68264
rect 0 65968 400 66024
rect 0 63728 400 63784
rect 0 61488 400 61544
rect 0 59248 400 59304
rect 0 57008 400 57064
rect 0 54768 400 54824
rect 0 52528 400 52584
rect 0 50288 400 50344
rect 0 48048 400 48104
rect 0 45808 400 45864
rect 0 43568 400 43624
rect 0 41328 400 41384
rect 0 39088 400 39144
rect 0 36848 400 36904
rect 0 34608 400 34664
rect 0 32368 400 32424
rect 0 30128 400 30184
rect 0 27888 400 27944
rect 0 25648 400 25704
rect 0 23408 400 23464
rect 0 21168 400 21224
rect 0 18928 400 18984
rect 0 16688 400 16744
rect 0 14448 400 14504
rect 0 12208 400 12264
rect 0 9968 400 10024
rect 0 7728 400 7784
rect 0 5488 400 5544
<< obsm3 >>
rect 9 294534 299367 299978
rect 430 294418 299367 294534
rect 9 292294 299367 294418
rect 430 292178 299367 292294
rect 9 290054 299367 292178
rect 430 289938 299367 290054
rect 9 287814 299367 289938
rect 430 287698 299367 287814
rect 9 285574 299367 287698
rect 430 285458 299367 285574
rect 9 283334 299367 285458
rect 430 283218 299367 283334
rect 9 281094 299367 283218
rect 430 280978 299367 281094
rect 9 278854 299367 280978
rect 430 278738 299367 278854
rect 9 276614 299367 278738
rect 430 276498 299367 276614
rect 9 274374 299367 276498
rect 430 274258 299367 274374
rect 9 272134 299367 274258
rect 430 272018 299367 272134
rect 9 269894 299367 272018
rect 430 269778 299367 269894
rect 9 267654 299367 269778
rect 430 267538 299367 267654
rect 9 265414 299367 267538
rect 430 265298 299367 265414
rect 9 263174 299367 265298
rect 430 263058 299367 263174
rect 9 260934 299367 263058
rect 430 260818 299367 260934
rect 9 258694 299367 260818
rect 430 258578 299367 258694
rect 9 256454 299367 258578
rect 430 256338 299367 256454
rect 9 254214 299367 256338
rect 430 254098 299367 254214
rect 9 251974 299367 254098
rect 430 251858 299367 251974
rect 9 249734 299367 251858
rect 430 249618 299367 249734
rect 9 247494 299367 249618
rect 430 247378 299367 247494
rect 9 245254 299367 247378
rect 430 245138 299367 245254
rect 9 243014 299367 245138
rect 430 242898 299367 243014
rect 9 240774 299367 242898
rect 430 240658 299367 240774
rect 9 238534 299367 240658
rect 430 238418 299367 238534
rect 9 236294 299367 238418
rect 430 236178 299367 236294
rect 9 234054 299367 236178
rect 430 233938 299367 234054
rect 9 231814 299367 233938
rect 430 231698 299367 231814
rect 9 229574 299367 231698
rect 430 229458 299367 229574
rect 9 227334 299367 229458
rect 430 227218 299367 227334
rect 9 225094 299367 227218
rect 430 224978 299367 225094
rect 9 222854 299367 224978
rect 430 222738 299367 222854
rect 9 220614 299367 222738
rect 430 220498 299367 220614
rect 9 218374 299367 220498
rect 430 218258 299367 218374
rect 9 216134 299367 218258
rect 430 216018 299367 216134
rect 9 213894 299367 216018
rect 430 213778 299367 213894
rect 9 211654 299367 213778
rect 430 211538 299367 211654
rect 9 209414 299367 211538
rect 430 209298 299367 209414
rect 9 207174 299367 209298
rect 430 207058 299367 207174
rect 9 204934 299367 207058
rect 430 204818 299367 204934
rect 9 202694 299367 204818
rect 430 202578 299367 202694
rect 9 200454 299367 202578
rect 430 200338 299367 200454
rect 9 198214 299367 200338
rect 430 198098 299367 198214
rect 9 195974 299367 198098
rect 430 195858 299367 195974
rect 9 193734 299367 195858
rect 430 193618 299367 193734
rect 9 191494 299367 193618
rect 430 191378 299367 191494
rect 9 189254 299367 191378
rect 430 189138 299367 189254
rect 9 187014 299367 189138
rect 430 186898 299367 187014
rect 9 184774 299367 186898
rect 430 184658 299367 184774
rect 9 182534 299367 184658
rect 430 182418 299367 182534
rect 9 180294 299367 182418
rect 430 180178 299367 180294
rect 9 178054 299367 180178
rect 430 177938 299367 178054
rect 9 175814 299367 177938
rect 430 175698 299367 175814
rect 9 173574 299367 175698
rect 430 173458 299367 173574
rect 9 171334 299367 173458
rect 430 171218 299367 171334
rect 9 169094 299367 171218
rect 430 168978 299367 169094
rect 9 166854 299367 168978
rect 430 166738 299367 166854
rect 9 164614 299367 166738
rect 430 164498 299367 164614
rect 9 162374 299367 164498
rect 430 162258 299367 162374
rect 9 160134 299367 162258
rect 430 160018 299367 160134
rect 9 157894 299367 160018
rect 430 157778 299367 157894
rect 9 155654 299367 157778
rect 430 155538 299367 155654
rect 9 153414 299367 155538
rect 430 153298 299367 153414
rect 9 151174 299367 153298
rect 430 151058 299367 151174
rect 9 148934 299367 151058
rect 430 148818 299367 148934
rect 9 146694 299367 148818
rect 430 146578 299367 146694
rect 9 144454 299367 146578
rect 430 144338 299367 144454
rect 9 142214 299367 144338
rect 430 142098 299367 142214
rect 9 139974 299367 142098
rect 430 139858 299367 139974
rect 9 137734 299367 139858
rect 430 137618 299367 137734
rect 9 135494 299367 137618
rect 430 135378 299367 135494
rect 9 133254 299367 135378
rect 430 133138 299367 133254
rect 9 131014 299367 133138
rect 430 130898 299367 131014
rect 9 128774 299367 130898
rect 430 128658 299367 128774
rect 9 126534 299367 128658
rect 430 126418 299367 126534
rect 9 124294 299367 126418
rect 430 124178 299367 124294
rect 9 122054 299367 124178
rect 430 121938 299367 122054
rect 9 119814 299367 121938
rect 430 119698 299367 119814
rect 9 117574 299367 119698
rect 430 117458 299367 117574
rect 9 115334 299367 117458
rect 430 115218 299367 115334
rect 9 113094 299367 115218
rect 430 112978 299367 113094
rect 9 110854 299367 112978
rect 430 110738 299367 110854
rect 9 108614 299367 110738
rect 430 108498 299367 108614
rect 9 106374 299367 108498
rect 430 106258 299367 106374
rect 9 104134 299367 106258
rect 430 104018 299367 104134
rect 9 101894 299367 104018
rect 430 101778 299367 101894
rect 9 99654 299367 101778
rect 430 99538 299367 99654
rect 9 97414 299367 99538
rect 430 97298 299367 97414
rect 9 95174 299367 97298
rect 430 95058 299367 95174
rect 9 92934 299367 95058
rect 430 92818 299367 92934
rect 9 90694 299367 92818
rect 430 90578 299367 90694
rect 9 88454 299367 90578
rect 430 88338 299367 88454
rect 9 86214 299367 88338
rect 430 86098 299367 86214
rect 9 83974 299367 86098
rect 430 83858 299367 83974
rect 9 81734 299367 83858
rect 430 81618 299367 81734
rect 9 79494 299367 81618
rect 430 79378 299367 79494
rect 9 77254 299367 79378
rect 430 77138 299367 77254
rect 9 75014 299367 77138
rect 430 74898 299367 75014
rect 9 72774 299367 74898
rect 430 72658 299367 72774
rect 9 70534 299367 72658
rect 430 70418 299367 70534
rect 9 68294 299367 70418
rect 430 68178 299367 68294
rect 9 66054 299367 68178
rect 430 65938 299367 66054
rect 9 63814 299367 65938
rect 430 63698 299367 63814
rect 9 61574 299367 63698
rect 430 61458 299367 61574
rect 9 59334 299367 61458
rect 430 59218 299367 59334
rect 9 57094 299367 59218
rect 430 56978 299367 57094
rect 9 54854 299367 56978
rect 430 54738 299367 54854
rect 9 52614 299367 54738
rect 430 52498 299367 52614
rect 9 50374 299367 52498
rect 430 50258 299367 50374
rect 9 48134 299367 50258
rect 430 48018 299367 48134
rect 9 45894 299367 48018
rect 430 45778 299367 45894
rect 9 43654 299367 45778
rect 430 43538 299367 43654
rect 9 41414 299367 43538
rect 430 41298 299367 41414
rect 9 39174 299367 41298
rect 430 39058 299367 39174
rect 9 36934 299367 39058
rect 430 36818 299367 36934
rect 9 34694 299367 36818
rect 430 34578 299367 34694
rect 9 32454 299367 34578
rect 430 32338 299367 32454
rect 9 30214 299367 32338
rect 430 30098 299367 30214
rect 9 27974 299367 30098
rect 430 27858 299367 27974
rect 9 25734 299367 27858
rect 430 25618 299367 25734
rect 9 23494 299367 25618
rect 430 23378 299367 23494
rect 9 21254 299367 23378
rect 430 21138 299367 21254
rect 9 19014 299367 21138
rect 430 18898 299367 19014
rect 9 16774 299367 18898
rect 430 16658 299367 16774
rect 9 14534 299367 16658
rect 430 14418 299367 14534
rect 9 12294 299367 14418
rect 430 12178 299367 12294
rect 9 10054 299367 12178
rect 430 9938 299367 10054
rect 9 7814 299367 9938
rect 430 7698 299367 7814
rect 9 5574 299367 7698
rect 430 5458 299367 5574
rect 9 14 299367 5458
<< metal4 >>
rect 2224 1538 2384 298342
rect 9904 1538 10064 298342
rect 17584 1538 17744 298342
rect 25264 1538 25424 298342
rect 32944 1538 33104 298342
rect 40624 1538 40784 298342
rect 48304 1538 48464 298342
rect 55984 1538 56144 298342
rect 63664 1538 63824 298342
rect 71344 1538 71504 298342
rect 79024 1538 79184 298342
rect 86704 1538 86864 298342
rect 94384 1538 94544 298342
rect 102064 1538 102224 298342
rect 109744 1538 109904 298342
rect 117424 1538 117584 298342
rect 125104 1538 125264 298342
rect 132784 1538 132944 298342
rect 140464 1538 140624 298342
rect 148144 1538 148304 298342
rect 155824 1538 155984 298342
rect 163504 1538 163664 298342
rect 171184 1538 171344 298342
rect 178864 1538 179024 298342
rect 186544 1538 186704 298342
rect 194224 1538 194384 298342
rect 201904 1538 202064 298342
rect 209584 1538 209744 298342
rect 217264 1538 217424 298342
rect 224944 1538 225104 298342
rect 232624 1538 232784 298342
rect 240304 1538 240464 298342
rect 247984 1538 248144 298342
rect 255664 1538 255824 298342
rect 263344 1538 263504 298342
rect 271024 1538 271184 298342
rect 278704 1538 278864 298342
rect 286384 1538 286544 298342
rect 294064 1538 294224 298342
<< obsm4 >>
rect 798 298372 298970 299983
rect 798 1508 2194 298372
rect 2414 1508 9874 298372
rect 10094 1508 17554 298372
rect 17774 1508 25234 298372
rect 25454 1508 32914 298372
rect 33134 1508 40594 298372
rect 40814 1508 48274 298372
rect 48494 1508 55954 298372
rect 56174 1508 63634 298372
rect 63854 1508 71314 298372
rect 71534 1508 78994 298372
rect 79214 1508 86674 298372
rect 86894 1508 94354 298372
rect 94574 1508 102034 298372
rect 102254 1508 109714 298372
rect 109934 1508 117394 298372
rect 117614 1508 125074 298372
rect 125294 1508 132754 298372
rect 132974 1508 140434 298372
rect 140654 1508 148114 298372
rect 148334 1508 155794 298372
rect 156014 1508 163474 298372
rect 163694 1508 171154 298372
rect 171374 1508 178834 298372
rect 179054 1508 186514 298372
rect 186734 1508 194194 298372
rect 194414 1508 201874 298372
rect 202094 1508 209554 298372
rect 209774 1508 217234 298372
rect 217454 1508 224914 298372
rect 225134 1508 232594 298372
rect 232814 1508 240274 298372
rect 240494 1508 247954 298372
rect 248174 1508 255634 298372
rect 255854 1508 263314 298372
rect 263534 1508 270994 298372
rect 271214 1508 278674 298372
rect 278894 1508 286354 298372
rect 286574 1508 294034 298372
rect 294254 1508 298970 298372
rect 798 9 298970 1508
<< labels >>
rlabel metal2 s 46928 299600 46984 300000 6 IN_DCT_data[0]
port 1 nsew signal input
rlabel metal2 s 24528 299600 24584 300000 6 IN_DCT_data[10]
port 2 nsew signal input
rlabel metal2 s 22288 299600 22344 300000 6 IN_DCT_data[11]
port 3 nsew signal input
rlabel metal2 s 20048 299600 20104 300000 6 IN_DCT_data[12]
port 4 nsew signal input
rlabel metal2 s 17808 299600 17864 300000 6 IN_DCT_data[13]
port 5 nsew signal input
rlabel metal2 s 15568 299600 15624 300000 6 IN_DCT_data[14]
port 6 nsew signal input
rlabel metal2 s 13328 299600 13384 300000 6 IN_DCT_data[15]
port 7 nsew signal input
rlabel metal2 s 11088 299600 11144 300000 6 IN_DCT_data[16]
port 8 nsew signal input
rlabel metal2 s 8848 299600 8904 300000 6 IN_DCT_data[17]
port 9 nsew signal input
rlabel metal2 s 6608 299600 6664 300000 6 IN_DCT_data[18]
port 10 nsew signal input
rlabel metal2 s 4368 299600 4424 300000 6 IN_DCT_data[19]
port 11 nsew signal input
rlabel metal2 s 44688 299600 44744 300000 6 IN_DCT_data[1]
port 12 nsew signal input
rlabel metal2 s 2128 299600 2184 300000 6 IN_DCT_data[20]
port 13 nsew signal input
rlabel metal2 s 42448 299600 42504 300000 6 IN_DCT_data[2]
port 14 nsew signal input
rlabel metal2 s 40208 299600 40264 300000 6 IN_DCT_data[3]
port 15 nsew signal input
rlabel metal2 s 37968 299600 38024 300000 6 IN_DCT_data[4]
port 16 nsew signal input
rlabel metal2 s 35728 299600 35784 300000 6 IN_DCT_data[5]
port 17 nsew signal input
rlabel metal2 s 33488 299600 33544 300000 6 IN_DCT_data[6]
port 18 nsew signal input
rlabel metal2 s 31248 299600 31304 300000 6 IN_DCT_data[7]
port 19 nsew signal input
rlabel metal2 s 29008 299600 29064 300000 6 IN_DCT_data[8]
port 20 nsew signal input
rlabel metal2 s 26768 299600 26824 300000 6 IN_DCT_data[9]
port 21 nsew signal input
rlabel metal2 s 190288 299600 190344 300000 6 IN_DC_data[0]
port 22 nsew signal input
rlabel metal2 s 167888 299600 167944 300000 6 IN_DC_data[10]
port 23 nsew signal input
rlabel metal2 s 165648 299600 165704 300000 6 IN_DC_data[11]
port 24 nsew signal input
rlabel metal2 s 163408 299600 163464 300000 6 IN_DC_data[12]
port 25 nsew signal input
rlabel metal2 s 161168 299600 161224 300000 6 IN_DC_data[13]
port 26 nsew signal input
rlabel metal2 s 158928 299600 158984 300000 6 IN_DC_data[14]
port 27 nsew signal input
rlabel metal2 s 156688 299600 156744 300000 6 IN_DC_data[15]
port 28 nsew signal input
rlabel metal2 s 154448 299600 154504 300000 6 IN_DC_data[16]
port 29 nsew signal input
rlabel metal2 s 152208 299600 152264 300000 6 IN_DC_data[17]
port 30 nsew signal input
rlabel metal2 s 149968 299600 150024 300000 6 IN_DC_data[18]
port 31 nsew signal input
rlabel metal2 s 147728 299600 147784 300000 6 IN_DC_data[19]
port 32 nsew signal input
rlabel metal2 s 188048 299600 188104 300000 6 IN_DC_data[1]
port 33 nsew signal input
rlabel metal2 s 145488 299600 145544 300000 6 IN_DC_data[20]
port 34 nsew signal input
rlabel metal2 s 143248 299600 143304 300000 6 IN_DC_data[21]
port 35 nsew signal input
rlabel metal2 s 141008 299600 141064 300000 6 IN_DC_data[22]
port 36 nsew signal input
rlabel metal2 s 138768 299600 138824 300000 6 IN_DC_data[23]
port 37 nsew signal input
rlabel metal2 s 136528 299600 136584 300000 6 IN_DC_data[24]
port 38 nsew signal input
rlabel metal2 s 134288 299600 134344 300000 6 IN_DC_data[25]
port 39 nsew signal input
rlabel metal2 s 132048 299600 132104 300000 6 IN_DC_data[26]
port 40 nsew signal input
rlabel metal2 s 129808 299600 129864 300000 6 IN_DC_data[27]
port 41 nsew signal input
rlabel metal2 s 127568 299600 127624 300000 6 IN_DC_data[28]
port 42 nsew signal input
rlabel metal2 s 125328 299600 125384 300000 6 IN_DC_data[29]
port 43 nsew signal input
rlabel metal2 s 185808 299600 185864 300000 6 IN_DC_data[2]
port 44 nsew signal input
rlabel metal2 s 123088 299600 123144 300000 6 IN_DC_data[30]
port 45 nsew signal input
rlabel metal2 s 120848 299600 120904 300000 6 IN_DC_data[31]
port 46 nsew signal input
rlabel metal2 s 183568 299600 183624 300000 6 IN_DC_data[3]
port 47 nsew signal input
rlabel metal2 s 181328 299600 181384 300000 6 IN_DC_data[4]
port 48 nsew signal input
rlabel metal2 s 179088 299600 179144 300000 6 IN_DC_data[5]
port 49 nsew signal input
rlabel metal2 s 176848 299600 176904 300000 6 IN_DC_data[6]
port 50 nsew signal input
rlabel metal2 s 174608 299600 174664 300000 6 IN_DC_data[7]
port 51 nsew signal input
rlabel metal2 s 172368 299600 172424 300000 6 IN_DC_data[8]
port 52 nsew signal input
rlabel metal2 s 170128 299600 170184 300000 6 IN_DC_data[9]
port 53 nsew signal input
rlabel metal3 s 0 50288 400 50344 6 IN_ICT_data[0]
port 54 nsew signal input
rlabel metal3 s 0 27888 400 27944 6 IN_ICT_data[10]
port 55 nsew signal input
rlabel metal3 s 0 25648 400 25704 6 IN_ICT_data[11]
port 56 nsew signal input
rlabel metal3 s 0 23408 400 23464 6 IN_ICT_data[12]
port 57 nsew signal input
rlabel metal3 s 0 21168 400 21224 6 IN_ICT_data[13]
port 58 nsew signal input
rlabel metal3 s 0 18928 400 18984 6 IN_ICT_data[14]
port 59 nsew signal input
rlabel metal3 s 0 16688 400 16744 6 IN_ICT_data[15]
port 60 nsew signal input
rlabel metal3 s 0 14448 400 14504 6 IN_ICT_data[16]
port 61 nsew signal input
rlabel metal3 s 0 12208 400 12264 6 IN_ICT_data[17]
port 62 nsew signal input
rlabel metal3 s 0 9968 400 10024 6 IN_ICT_data[18]
port 63 nsew signal input
rlabel metal3 s 0 7728 400 7784 6 IN_ICT_data[19]
port 64 nsew signal input
rlabel metal3 s 0 48048 400 48104 6 IN_ICT_data[1]
port 65 nsew signal input
rlabel metal3 s 0 5488 400 5544 6 IN_ICT_data[20]
port 66 nsew signal input
rlabel metal3 s 0 45808 400 45864 6 IN_ICT_data[2]
port 67 nsew signal input
rlabel metal3 s 0 43568 400 43624 6 IN_ICT_data[3]
port 68 nsew signal input
rlabel metal3 s 0 41328 400 41384 6 IN_ICT_data[4]
port 69 nsew signal input
rlabel metal3 s 0 39088 400 39144 6 IN_ICT_data[5]
port 70 nsew signal input
rlabel metal3 s 0 36848 400 36904 6 IN_ICT_data[6]
port 71 nsew signal input
rlabel metal3 s 0 34608 400 34664 6 IN_ICT_data[7]
port 72 nsew signal input
rlabel metal3 s 0 32368 400 32424 6 IN_ICT_data[8]
port 73 nsew signal input
rlabel metal3 s 0 30128 400 30184 6 IN_ICT_data[9]
port 74 nsew signal input
rlabel metal3 s 0 193648 400 193704 6 IN_IC_data[0]
port 75 nsew signal input
rlabel metal3 s 0 171248 400 171304 6 IN_IC_data[10]
port 76 nsew signal input
rlabel metal3 s 0 169008 400 169064 6 IN_IC_data[11]
port 77 nsew signal input
rlabel metal3 s 0 166768 400 166824 6 IN_IC_data[12]
port 78 nsew signal input
rlabel metal3 s 0 164528 400 164584 6 IN_IC_data[13]
port 79 nsew signal input
rlabel metal3 s 0 162288 400 162344 6 IN_IC_data[14]
port 80 nsew signal input
rlabel metal3 s 0 160048 400 160104 6 IN_IC_data[15]
port 81 nsew signal input
rlabel metal3 s 0 157808 400 157864 6 IN_IC_data[16]
port 82 nsew signal input
rlabel metal3 s 0 155568 400 155624 6 IN_IC_data[17]
port 83 nsew signal input
rlabel metal3 s 0 153328 400 153384 6 IN_IC_data[18]
port 84 nsew signal input
rlabel metal3 s 0 151088 400 151144 6 IN_IC_data[19]
port 85 nsew signal input
rlabel metal3 s 0 191408 400 191464 6 IN_IC_data[1]
port 86 nsew signal input
rlabel metal3 s 0 148848 400 148904 6 IN_IC_data[20]
port 87 nsew signal input
rlabel metal3 s 0 146608 400 146664 6 IN_IC_data[21]
port 88 nsew signal input
rlabel metal3 s 0 144368 400 144424 6 IN_IC_data[22]
port 89 nsew signal input
rlabel metal3 s 0 142128 400 142184 6 IN_IC_data[23]
port 90 nsew signal input
rlabel metal3 s 0 139888 400 139944 6 IN_IC_data[24]
port 91 nsew signal input
rlabel metal3 s 0 137648 400 137704 6 IN_IC_data[25]
port 92 nsew signal input
rlabel metal3 s 0 135408 400 135464 6 IN_IC_data[26]
port 93 nsew signal input
rlabel metal3 s 0 133168 400 133224 6 IN_IC_data[27]
port 94 nsew signal input
rlabel metal3 s 0 130928 400 130984 6 IN_IC_data[28]
port 95 nsew signal input
rlabel metal3 s 0 128688 400 128744 6 IN_IC_data[29]
port 96 nsew signal input
rlabel metal3 s 0 189168 400 189224 6 IN_IC_data[2]
port 97 nsew signal input
rlabel metal3 s 0 126448 400 126504 6 IN_IC_data[30]
port 98 nsew signal input
rlabel metal3 s 0 124208 400 124264 6 IN_IC_data[31]
port 99 nsew signal input
rlabel metal3 s 0 186928 400 186984 6 IN_IC_data[3]
port 100 nsew signal input
rlabel metal3 s 0 184688 400 184744 6 IN_IC_data[4]
port 101 nsew signal input
rlabel metal3 s 0 182448 400 182504 6 IN_IC_data[5]
port 102 nsew signal input
rlabel metal3 s 0 180208 400 180264 6 IN_IC_data[6]
port 103 nsew signal input
rlabel metal3 s 0 177968 400 178024 6 IN_IC_data[7]
port 104 nsew signal input
rlabel metal3 s 0 175728 400 175784 6 IN_IC_data[8]
port 105 nsew signal input
rlabel metal3 s 0 173488 400 173544 6 IN_IC_data[9]
port 106 nsew signal input
rlabel metal2 s 111888 299600 111944 300000 6 OUT_DCT_addr[0]
port 107 nsew signal output
rlabel metal2 s 107408 299600 107464 300000 6 OUT_DCT_addr[1]
port 108 nsew signal output
rlabel metal2 s 102928 299600 102984 300000 6 OUT_DCT_addr[2]
port 109 nsew signal output
rlabel metal2 s 98448 299600 98504 300000 6 OUT_DCT_addr[3]
port 110 nsew signal output
rlabel metal2 s 93968 299600 94024 300000 6 OUT_DCT_addr[4]
port 111 nsew signal output
rlabel metal2 s 89488 299600 89544 300000 6 OUT_DCT_addr[5]
port 112 nsew signal output
rlabel metal2 s 85008 299600 85064 300000 6 OUT_DCT_addr[6]
port 113 nsew signal output
rlabel metal2 s 80528 299600 80584 300000 6 OUT_DCT_addr[7]
port 114 nsew signal output
rlabel metal2 s 118608 299600 118664 300000 6 OUT_DCT_ce
port 115 nsew signal output
rlabel metal2 s 109648 299600 109704 300000 6 OUT_DCT_data[0]
port 116 nsew signal output
rlabel metal2 s 71568 299600 71624 300000 6 OUT_DCT_data[10]
port 117 nsew signal output
rlabel metal2 s 69328 299600 69384 300000 6 OUT_DCT_data[11]
port 118 nsew signal output
rlabel metal2 s 67088 299600 67144 300000 6 OUT_DCT_data[12]
port 119 nsew signal output
rlabel metal2 s 64848 299600 64904 300000 6 OUT_DCT_data[13]
port 120 nsew signal output
rlabel metal2 s 62608 299600 62664 300000 6 OUT_DCT_data[14]
port 121 nsew signal output
rlabel metal2 s 60368 299600 60424 300000 6 OUT_DCT_data[15]
port 122 nsew signal output
rlabel metal2 s 58128 299600 58184 300000 6 OUT_DCT_data[16]
port 123 nsew signal output
rlabel metal2 s 55888 299600 55944 300000 6 OUT_DCT_data[17]
port 124 nsew signal output
rlabel metal2 s 53648 299600 53704 300000 6 OUT_DCT_data[18]
port 125 nsew signal output
rlabel metal2 s 51408 299600 51464 300000 6 OUT_DCT_data[19]
port 126 nsew signal output
rlabel metal2 s 105168 299600 105224 300000 6 OUT_DCT_data[1]
port 127 nsew signal output
rlabel metal2 s 49168 299600 49224 300000 6 OUT_DCT_data[20]
port 128 nsew signal output
rlabel metal2 s 100688 299600 100744 300000 6 OUT_DCT_data[2]
port 129 nsew signal output
rlabel metal2 s 96208 299600 96264 300000 6 OUT_DCT_data[3]
port 130 nsew signal output
rlabel metal2 s 91728 299600 91784 300000 6 OUT_DCT_data[4]
port 131 nsew signal output
rlabel metal2 s 87248 299600 87304 300000 6 OUT_DCT_data[5]
port 132 nsew signal output
rlabel metal2 s 82768 299600 82824 300000 6 OUT_DCT_data[6]
port 133 nsew signal output
rlabel metal2 s 78288 299600 78344 300000 6 OUT_DCT_data[7]
port 134 nsew signal output
rlabel metal2 s 76048 299600 76104 300000 6 OUT_DCT_data[8]
port 135 nsew signal output
rlabel metal2 s 73808 299600 73864 300000 6 OUT_DCT_data[9]
port 136 nsew signal output
rlabel metal2 s 116368 299600 116424 300000 6 OUT_DCT_we
port 137 nsew signal output
rlabel metal2 s 114128 299600 114184 300000 6 OUT_DCT_wm
port 138 nsew signal output
rlabel metal2 s 293328 299600 293384 300000 6 OUT_DC_addr[0]
port 139 nsew signal output
rlabel metal2 s 286608 299600 286664 300000 6 OUT_DC_addr[1]
port 140 nsew signal output
rlabel metal2 s 279888 299600 279944 300000 6 OUT_DC_addr[2]
port 141 nsew signal output
rlabel metal2 s 273168 299600 273224 300000 6 OUT_DC_addr[3]
port 142 nsew signal output
rlabel metal2 s 266448 299600 266504 300000 6 OUT_DC_addr[4]
port 143 nsew signal output
rlabel metal2 s 261968 299600 262024 300000 6 OUT_DC_addr[5]
port 144 nsew signal output
rlabel metal2 s 257488 299600 257544 300000 6 OUT_DC_addr[6]
port 145 nsew signal output
rlabel metal2 s 253008 299600 253064 300000 6 OUT_DC_addr[7]
port 146 nsew signal output
rlabel metal2 s 248528 299600 248584 300000 6 OUT_DC_addr[8]
port 147 nsew signal output
rlabel metal2 s 244048 299600 244104 300000 6 OUT_DC_addr[9]
port 148 nsew signal output
rlabel metal2 s 297808 299600 297864 300000 6 OUT_DC_ce
port 149 nsew signal output
rlabel metal2 s 291088 299600 291144 300000 6 OUT_DC_data[0]
port 150 nsew signal output
rlabel metal2 s 239568 299600 239624 300000 6 OUT_DC_data[10]
port 151 nsew signal output
rlabel metal2 s 237328 299600 237384 300000 6 OUT_DC_data[11]
port 152 nsew signal output
rlabel metal2 s 235088 299600 235144 300000 6 OUT_DC_data[12]
port 153 nsew signal output
rlabel metal2 s 232848 299600 232904 300000 6 OUT_DC_data[13]
port 154 nsew signal output
rlabel metal2 s 230608 299600 230664 300000 6 OUT_DC_data[14]
port 155 nsew signal output
rlabel metal2 s 228368 299600 228424 300000 6 OUT_DC_data[15]
port 156 nsew signal output
rlabel metal2 s 226128 299600 226184 300000 6 OUT_DC_data[16]
port 157 nsew signal output
rlabel metal2 s 223888 299600 223944 300000 6 OUT_DC_data[17]
port 158 nsew signal output
rlabel metal2 s 221648 299600 221704 300000 6 OUT_DC_data[18]
port 159 nsew signal output
rlabel metal2 s 219408 299600 219464 300000 6 OUT_DC_data[19]
port 160 nsew signal output
rlabel metal2 s 284368 299600 284424 300000 6 OUT_DC_data[1]
port 161 nsew signal output
rlabel metal2 s 217168 299600 217224 300000 6 OUT_DC_data[20]
port 162 nsew signal output
rlabel metal2 s 214928 299600 214984 300000 6 OUT_DC_data[21]
port 163 nsew signal output
rlabel metal2 s 212688 299600 212744 300000 6 OUT_DC_data[22]
port 164 nsew signal output
rlabel metal2 s 210448 299600 210504 300000 6 OUT_DC_data[23]
port 165 nsew signal output
rlabel metal2 s 208208 299600 208264 300000 6 OUT_DC_data[24]
port 166 nsew signal output
rlabel metal2 s 205968 299600 206024 300000 6 OUT_DC_data[25]
port 167 nsew signal output
rlabel metal2 s 203728 299600 203784 300000 6 OUT_DC_data[26]
port 168 nsew signal output
rlabel metal2 s 201488 299600 201544 300000 6 OUT_DC_data[27]
port 169 nsew signal output
rlabel metal2 s 199248 299600 199304 300000 6 OUT_DC_data[28]
port 170 nsew signal output
rlabel metal2 s 197008 299600 197064 300000 6 OUT_DC_data[29]
port 171 nsew signal output
rlabel metal2 s 277648 299600 277704 300000 6 OUT_DC_data[2]
port 172 nsew signal output
rlabel metal2 s 194768 299600 194824 300000 6 OUT_DC_data[30]
port 173 nsew signal output
rlabel metal2 s 192528 299600 192584 300000 6 OUT_DC_data[31]
port 174 nsew signal output
rlabel metal2 s 270928 299600 270984 300000 6 OUT_DC_data[3]
port 175 nsew signal output
rlabel metal2 s 264208 299600 264264 300000 6 OUT_DC_data[4]
port 176 nsew signal output
rlabel metal2 s 259728 299600 259784 300000 6 OUT_DC_data[5]
port 177 nsew signal output
rlabel metal2 s 255248 299600 255304 300000 6 OUT_DC_data[6]
port 178 nsew signal output
rlabel metal2 s 250768 299600 250824 300000 6 OUT_DC_data[7]
port 179 nsew signal output
rlabel metal2 s 246288 299600 246344 300000 6 OUT_DC_data[8]
port 180 nsew signal output
rlabel metal2 s 241808 299600 241864 300000 6 OUT_DC_data[9]
port 181 nsew signal output
rlabel metal2 s 295568 299600 295624 300000 6 OUT_DC_we
port 182 nsew signal output
rlabel metal2 s 288848 299600 288904 300000 6 OUT_DC_wm[0]
port 183 nsew signal output
rlabel metal2 s 282128 299600 282184 300000 6 OUT_DC_wm[1]
port 184 nsew signal output
rlabel metal2 s 275408 299600 275464 300000 6 OUT_DC_wm[2]
port 185 nsew signal output
rlabel metal2 s 268688 299600 268744 300000 6 OUT_DC_wm[3]
port 186 nsew signal output
rlabel metal3 s 0 115248 400 115304 6 OUT_ICT_addr[0]
port 187 nsew signal output
rlabel metal3 s 0 110768 400 110824 6 OUT_ICT_addr[1]
port 188 nsew signal output
rlabel metal3 s 0 106288 400 106344 6 OUT_ICT_addr[2]
port 189 nsew signal output
rlabel metal3 s 0 101808 400 101864 6 OUT_ICT_addr[3]
port 190 nsew signal output
rlabel metal3 s 0 97328 400 97384 6 OUT_ICT_addr[4]
port 191 nsew signal output
rlabel metal3 s 0 92848 400 92904 6 OUT_ICT_addr[5]
port 192 nsew signal output
rlabel metal3 s 0 88368 400 88424 6 OUT_ICT_addr[6]
port 193 nsew signal output
rlabel metal3 s 0 83888 400 83944 6 OUT_ICT_addr[7]
port 194 nsew signal output
rlabel metal3 s 0 121968 400 122024 6 OUT_ICT_ce
port 195 nsew signal output
rlabel metal3 s 0 113008 400 113064 6 OUT_ICT_data[0]
port 196 nsew signal output
rlabel metal3 s 0 74928 400 74984 6 OUT_ICT_data[10]
port 197 nsew signal output
rlabel metal3 s 0 72688 400 72744 6 OUT_ICT_data[11]
port 198 nsew signal output
rlabel metal3 s 0 70448 400 70504 6 OUT_ICT_data[12]
port 199 nsew signal output
rlabel metal3 s 0 68208 400 68264 6 OUT_ICT_data[13]
port 200 nsew signal output
rlabel metal3 s 0 65968 400 66024 6 OUT_ICT_data[14]
port 201 nsew signal output
rlabel metal3 s 0 63728 400 63784 6 OUT_ICT_data[15]
port 202 nsew signal output
rlabel metal3 s 0 61488 400 61544 6 OUT_ICT_data[16]
port 203 nsew signal output
rlabel metal3 s 0 59248 400 59304 6 OUT_ICT_data[17]
port 204 nsew signal output
rlabel metal3 s 0 57008 400 57064 6 OUT_ICT_data[18]
port 205 nsew signal output
rlabel metal3 s 0 54768 400 54824 6 OUT_ICT_data[19]
port 206 nsew signal output
rlabel metal3 s 0 108528 400 108584 6 OUT_ICT_data[1]
port 207 nsew signal output
rlabel metal3 s 0 52528 400 52584 6 OUT_ICT_data[20]
port 208 nsew signal output
rlabel metal3 s 0 104048 400 104104 6 OUT_ICT_data[2]
port 209 nsew signal output
rlabel metal3 s 0 99568 400 99624 6 OUT_ICT_data[3]
port 210 nsew signal output
rlabel metal3 s 0 95088 400 95144 6 OUT_ICT_data[4]
port 211 nsew signal output
rlabel metal3 s 0 90608 400 90664 6 OUT_ICT_data[5]
port 212 nsew signal output
rlabel metal3 s 0 86128 400 86184 6 OUT_ICT_data[6]
port 213 nsew signal output
rlabel metal3 s 0 81648 400 81704 6 OUT_ICT_data[7]
port 214 nsew signal output
rlabel metal3 s 0 79408 400 79464 6 OUT_ICT_data[8]
port 215 nsew signal output
rlabel metal3 s 0 77168 400 77224 6 OUT_ICT_data[9]
port 216 nsew signal output
rlabel metal3 s 0 119728 400 119784 6 OUT_ICT_we
port 217 nsew signal output
rlabel metal3 s 0 117488 400 117544 6 OUT_ICT_wm
port 218 nsew signal output
rlabel metal3 s 0 287728 400 287784 6 OUT_IC_addr[0]
port 219 nsew signal output
rlabel metal3 s 0 283248 400 283304 6 OUT_IC_addr[1]
port 220 nsew signal output
rlabel metal3 s 0 278768 400 278824 6 OUT_IC_addr[2]
port 221 nsew signal output
rlabel metal3 s 0 274288 400 274344 6 OUT_IC_addr[3]
port 222 nsew signal output
rlabel metal3 s 0 269808 400 269864 6 OUT_IC_addr[4]
port 223 nsew signal output
rlabel metal3 s 0 265328 400 265384 6 OUT_IC_addr[5]
port 224 nsew signal output
rlabel metal3 s 0 260848 400 260904 6 OUT_IC_addr[6]
port 225 nsew signal output
rlabel metal3 s 0 256368 400 256424 6 OUT_IC_addr[7]
port 226 nsew signal output
rlabel metal3 s 0 251888 400 251944 6 OUT_IC_addr[8]
port 227 nsew signal output
rlabel metal3 s 0 247408 400 247464 6 OUT_IC_addr[9]
port 228 nsew signal output
rlabel metal3 s 0 294448 400 294504 6 OUT_IC_ce
port 229 nsew signal output
rlabel metal3 s 0 285488 400 285544 6 OUT_IC_data[0]
port 230 nsew signal output
rlabel metal3 s 0 242928 400 242984 6 OUT_IC_data[10]
port 231 nsew signal output
rlabel metal3 s 0 240688 400 240744 6 OUT_IC_data[11]
port 232 nsew signal output
rlabel metal3 s 0 238448 400 238504 6 OUT_IC_data[12]
port 233 nsew signal output
rlabel metal3 s 0 236208 400 236264 6 OUT_IC_data[13]
port 234 nsew signal output
rlabel metal3 s 0 233968 400 234024 6 OUT_IC_data[14]
port 235 nsew signal output
rlabel metal3 s 0 231728 400 231784 6 OUT_IC_data[15]
port 236 nsew signal output
rlabel metal3 s 0 229488 400 229544 6 OUT_IC_data[16]
port 237 nsew signal output
rlabel metal3 s 0 227248 400 227304 6 OUT_IC_data[17]
port 238 nsew signal output
rlabel metal3 s 0 225008 400 225064 6 OUT_IC_data[18]
port 239 nsew signal output
rlabel metal3 s 0 222768 400 222824 6 OUT_IC_data[19]
port 240 nsew signal output
rlabel metal3 s 0 281008 400 281064 6 OUT_IC_data[1]
port 241 nsew signal output
rlabel metal3 s 0 220528 400 220584 6 OUT_IC_data[20]
port 242 nsew signal output
rlabel metal3 s 0 218288 400 218344 6 OUT_IC_data[21]
port 243 nsew signal output
rlabel metal3 s 0 216048 400 216104 6 OUT_IC_data[22]
port 244 nsew signal output
rlabel metal3 s 0 213808 400 213864 6 OUT_IC_data[23]
port 245 nsew signal output
rlabel metal3 s 0 211568 400 211624 6 OUT_IC_data[24]
port 246 nsew signal output
rlabel metal3 s 0 209328 400 209384 6 OUT_IC_data[25]
port 247 nsew signal output
rlabel metal3 s 0 207088 400 207144 6 OUT_IC_data[26]
port 248 nsew signal output
rlabel metal3 s 0 204848 400 204904 6 OUT_IC_data[27]
port 249 nsew signal output
rlabel metal3 s 0 202608 400 202664 6 OUT_IC_data[28]
port 250 nsew signal output
rlabel metal3 s 0 200368 400 200424 6 OUT_IC_data[29]
port 251 nsew signal output
rlabel metal3 s 0 276528 400 276584 6 OUT_IC_data[2]
port 252 nsew signal output
rlabel metal3 s 0 198128 400 198184 6 OUT_IC_data[30]
port 253 nsew signal output
rlabel metal3 s 0 195888 400 195944 6 OUT_IC_data[31]
port 254 nsew signal output
rlabel metal3 s 0 272048 400 272104 6 OUT_IC_data[3]
port 255 nsew signal output
rlabel metal3 s 0 267568 400 267624 6 OUT_IC_data[4]
port 256 nsew signal output
rlabel metal3 s 0 263088 400 263144 6 OUT_IC_data[5]
port 257 nsew signal output
rlabel metal3 s 0 258608 400 258664 6 OUT_IC_data[6]
port 258 nsew signal output
rlabel metal3 s 0 254128 400 254184 6 OUT_IC_data[7]
port 259 nsew signal output
rlabel metal3 s 0 249648 400 249704 6 OUT_IC_data[8]
port 260 nsew signal output
rlabel metal3 s 0 245168 400 245224 6 OUT_IC_data[9]
port 261 nsew signal output
rlabel metal3 s 0 292208 400 292264 6 OUT_IC_we
port 262 nsew signal output
rlabel metal3 s 0 289968 400 290024 6 OUT_IC_wm
port 263 nsew signal output
rlabel metal2 s 226128 0 226184 400 6 OUT_dbgMemC[0]
port 264 nsew signal output
rlabel metal2 s 248528 0 248584 400 6 OUT_dbgMemC[10]
port 265 nsew signal output
rlabel metal2 s 250768 0 250824 400 6 OUT_dbgMemC[11]
port 266 nsew signal output
rlabel metal2 s 253008 0 253064 400 6 OUT_dbgMemC[12]
port 267 nsew signal output
rlabel metal2 s 255248 0 255304 400 6 OUT_dbgMemC[13]
port 268 nsew signal output
rlabel metal2 s 257488 0 257544 400 6 OUT_dbgMemC[14]
port 269 nsew signal output
rlabel metal2 s 259728 0 259784 400 6 OUT_dbgMemC[15]
port 270 nsew signal output
rlabel metal2 s 228368 0 228424 400 6 OUT_dbgMemC[1]
port 271 nsew signal output
rlabel metal2 s 230608 0 230664 400 6 OUT_dbgMemC[2]
port 272 nsew signal output
rlabel metal2 s 232848 0 232904 400 6 OUT_dbgMemC[3]
port 273 nsew signal output
rlabel metal2 s 235088 0 235144 400 6 OUT_dbgMemC[4]
port 274 nsew signal output
rlabel metal2 s 237328 0 237384 400 6 OUT_dbgMemC[5]
port 275 nsew signal output
rlabel metal2 s 239568 0 239624 400 6 OUT_dbgMemC[6]
port 276 nsew signal output
rlabel metal2 s 241808 0 241864 400 6 OUT_dbgMemC[7]
port 277 nsew signal output
rlabel metal2 s 244048 0 244104 400 6 OUT_dbgMemC[8]
port 278 nsew signal output
rlabel metal2 s 246288 0 246344 400 6 OUT_dbgMemC[9]
port 279 nsew signal output
rlabel metal2 s 225008 0 225064 400 6 OUT_dbg[0]
port 280 nsew signal output
rlabel metal2 s 247408 0 247464 400 6 OUT_dbg[10]
port 281 nsew signal output
rlabel metal2 s 249648 0 249704 400 6 OUT_dbg[11]
port 282 nsew signal output
rlabel metal2 s 251888 0 251944 400 6 OUT_dbg[12]
port 283 nsew signal output
rlabel metal2 s 254128 0 254184 400 6 OUT_dbg[13]
port 284 nsew signal output
rlabel metal2 s 256368 0 256424 400 6 OUT_dbg[14]
port 285 nsew signal output
rlabel metal2 s 258608 0 258664 400 6 OUT_dbg[15]
port 286 nsew signal output
rlabel metal2 s 260848 0 260904 400 6 OUT_dbg[16]
port 287 nsew signal output
rlabel metal2 s 261968 0 262024 400 6 OUT_dbg[17]
port 288 nsew signal output
rlabel metal2 s 263088 0 263144 400 6 OUT_dbg[18]
port 289 nsew signal output
rlabel metal2 s 264208 0 264264 400 6 OUT_dbg[19]
port 290 nsew signal output
rlabel metal2 s 227248 0 227304 400 6 OUT_dbg[1]
port 291 nsew signal output
rlabel metal2 s 265328 0 265384 400 6 OUT_dbg[20]
port 292 nsew signal output
rlabel metal2 s 266448 0 266504 400 6 OUT_dbg[21]
port 293 nsew signal output
rlabel metal2 s 267568 0 267624 400 6 OUT_dbg[22]
port 294 nsew signal output
rlabel metal2 s 268688 0 268744 400 6 OUT_dbg[23]
port 295 nsew signal output
rlabel metal2 s 269808 0 269864 400 6 OUT_dbg[24]
port 296 nsew signal output
rlabel metal2 s 270928 0 270984 400 6 OUT_dbg[25]
port 297 nsew signal output
rlabel metal2 s 272048 0 272104 400 6 OUT_dbg[26]
port 298 nsew signal output
rlabel metal2 s 273168 0 273224 400 6 OUT_dbg[27]
port 299 nsew signal output
rlabel metal2 s 274288 0 274344 400 6 OUT_dbg[28]
port 300 nsew signal output
rlabel metal2 s 275408 0 275464 400 6 OUT_dbg[29]
port 301 nsew signal output
rlabel metal2 s 229488 0 229544 400 6 OUT_dbg[2]
port 302 nsew signal output
rlabel metal2 s 276528 0 276584 400 6 OUT_dbg[30]
port 303 nsew signal output
rlabel metal2 s 277648 0 277704 400 6 OUT_dbg[31]
port 304 nsew signal output
rlabel metal2 s 278768 0 278824 400 6 OUT_dbg[32]
port 305 nsew signal output
rlabel metal2 s 279888 0 279944 400 6 OUT_dbg[33]
port 306 nsew signal output
rlabel metal2 s 281008 0 281064 400 6 OUT_dbg[34]
port 307 nsew signal output
rlabel metal2 s 282128 0 282184 400 6 OUT_dbg[35]
port 308 nsew signal output
rlabel metal2 s 283248 0 283304 400 6 OUT_dbg[36]
port 309 nsew signal output
rlabel metal2 s 284368 0 284424 400 6 OUT_dbg[37]
port 310 nsew signal output
rlabel metal2 s 285488 0 285544 400 6 OUT_dbg[38]
port 311 nsew signal output
rlabel metal2 s 286608 0 286664 400 6 OUT_dbg[39]
port 312 nsew signal output
rlabel metal2 s 231728 0 231784 400 6 OUT_dbg[3]
port 313 nsew signal output
rlabel metal2 s 233968 0 234024 400 6 OUT_dbg[4]
port 314 nsew signal output
rlabel metal2 s 236208 0 236264 400 6 OUT_dbg[5]
port 315 nsew signal output
rlabel metal2 s 238448 0 238504 400 6 OUT_dbg[6]
port 316 nsew signal output
rlabel metal2 s 240688 0 240744 400 6 OUT_dbg[7]
port 317 nsew signal output
rlabel metal2 s 242928 0 242984 400 6 OUT_dbg[8]
port 318 nsew signal output
rlabel metal2 s 245168 0 245224 400 6 OUT_dbg[9]
port 319 nsew signal output
rlabel metal2 s 222768 0 222824 400 6 OUT_powerOff
port 320 nsew signal output
rlabel metal2 s 223888 0 223944 400 6 OUT_reboot
port 321 nsew signal output
rlabel metal2 s 219408 0 219464 400 6 clk
port 322 nsew signal input
rlabel metal2 s 221648 0 221704 400 6 en
port 323 nsew signal input
rlabel metal2 s 220528 0 220584 400 6 rst
port 324 nsew signal input
rlabel metal2 s 33488 0 33544 400 6 s_axi_araddr[0]
port 325 nsew signal output
rlabel metal2 s 120848 0 120904 400 6 s_axi_araddr[10]
port 326 nsew signal output
rlabel metal2 s 125328 0 125384 400 6 s_axi_araddr[11]
port 327 nsew signal output
rlabel metal2 s 129808 0 129864 400 6 s_axi_araddr[12]
port 328 nsew signal output
rlabel metal2 s 134288 0 134344 400 6 s_axi_araddr[13]
port 329 nsew signal output
rlabel metal2 s 138768 0 138824 400 6 s_axi_araddr[14]
port 330 nsew signal output
rlabel metal2 s 143248 0 143304 400 6 s_axi_araddr[15]
port 331 nsew signal output
rlabel metal2 s 147728 0 147784 400 6 s_axi_araddr[16]
port 332 nsew signal output
rlabel metal2 s 152208 0 152264 400 6 s_axi_araddr[17]
port 333 nsew signal output
rlabel metal2 s 156688 0 156744 400 6 s_axi_araddr[18]
port 334 nsew signal output
rlabel metal2 s 161168 0 161224 400 6 s_axi_araddr[19]
port 335 nsew signal output
rlabel metal2 s 48048 0 48104 400 6 s_axi_araddr[1]
port 336 nsew signal output
rlabel metal2 s 165648 0 165704 400 6 s_axi_araddr[20]
port 337 nsew signal output
rlabel metal2 s 170128 0 170184 400 6 s_axi_araddr[21]
port 338 nsew signal output
rlabel metal2 s 174608 0 174664 400 6 s_axi_araddr[22]
port 339 nsew signal output
rlabel metal2 s 179088 0 179144 400 6 s_axi_araddr[23]
port 340 nsew signal output
rlabel metal2 s 183568 0 183624 400 6 s_axi_araddr[24]
port 341 nsew signal output
rlabel metal2 s 188048 0 188104 400 6 s_axi_araddr[25]
port 342 nsew signal output
rlabel metal2 s 192528 0 192584 400 6 s_axi_araddr[26]
port 343 nsew signal output
rlabel metal2 s 197008 0 197064 400 6 s_axi_araddr[27]
port 344 nsew signal output
rlabel metal2 s 201488 0 201544 400 6 s_axi_araddr[28]
port 345 nsew signal output
rlabel metal2 s 205968 0 206024 400 6 s_axi_araddr[29]
port 346 nsew signal output
rlabel metal2 s 62608 0 62664 400 6 s_axi_araddr[2]
port 347 nsew signal output
rlabel metal2 s 210448 0 210504 400 6 s_axi_araddr[30]
port 348 nsew signal output
rlabel metal2 s 214928 0 214984 400 6 s_axi_araddr[31]
port 349 nsew signal output
rlabel metal2 s 74928 0 74984 400 6 s_axi_araddr[3]
port 350 nsew signal output
rlabel metal2 s 85008 0 85064 400 6 s_axi_araddr[4]
port 351 nsew signal output
rlabel metal2 s 91728 0 91784 400 6 s_axi_araddr[5]
port 352 nsew signal output
rlabel metal2 s 98448 0 98504 400 6 s_axi_araddr[6]
port 353 nsew signal output
rlabel metal2 s 105168 0 105224 400 6 s_axi_araddr[7]
port 354 nsew signal output
rlabel metal2 s 111888 0 111944 400 6 s_axi_araddr[8]
port 355 nsew signal output
rlabel metal2 s 116368 0 116424 400 6 s_axi_araddr[9]
port 356 nsew signal output
rlabel metal2 s 34608 0 34664 400 6 s_axi_arburst[0]
port 357 nsew signal output
rlabel metal2 s 49168 0 49224 400 6 s_axi_arburst[1]
port 358 nsew signal output
rlabel metal2 s 35728 0 35784 400 6 s_axi_arcache[0]
port 359 nsew signal output
rlabel metal2 s 50288 0 50344 400 6 s_axi_arcache[1]
port 360 nsew signal output
rlabel metal2 s 63728 0 63784 400 6 s_axi_arcache[2]
port 361 nsew signal output
rlabel metal2 s 76048 0 76104 400 6 s_axi_arcache[3]
port 362 nsew signal output
rlabel metal2 s 13328 0 13384 400 6 s_axi_arid
port 363 nsew signal output
rlabel metal2 s 36848 0 36904 400 6 s_axi_arlen[0]
port 364 nsew signal output
rlabel metal2 s 51408 0 51464 400 6 s_axi_arlen[1]
port 365 nsew signal output
rlabel metal2 s 64848 0 64904 400 6 s_axi_arlen[2]
port 366 nsew signal output
rlabel metal2 s 77168 0 77224 400 6 s_axi_arlen[3]
port 367 nsew signal output
rlabel metal2 s 86128 0 86184 400 6 s_axi_arlen[4]
port 368 nsew signal output
rlabel metal2 s 92848 0 92904 400 6 s_axi_arlen[5]
port 369 nsew signal output
rlabel metal2 s 99568 0 99624 400 6 s_axi_arlen[6]
port 370 nsew signal output
rlabel metal2 s 106288 0 106344 400 6 s_axi_arlen[7]
port 371 nsew signal output
rlabel metal2 s 14448 0 14504 400 6 s_axi_arlock
port 372 nsew signal output
rlabel metal2 s 15568 0 15624 400 6 s_axi_arready
port 373 nsew signal input
rlabel metal2 s 37968 0 38024 400 6 s_axi_arsize[0]
port 374 nsew signal output
rlabel metal2 s 52528 0 52584 400 6 s_axi_arsize[1]
port 375 nsew signal output
rlabel metal2 s 65968 0 66024 400 6 s_axi_arsize[2]
port 376 nsew signal output
rlabel metal2 s 16688 0 16744 400 6 s_axi_arvalid
port 377 nsew signal output
rlabel metal2 s 39088 0 39144 400 6 s_axi_awaddr[0]
port 378 nsew signal output
rlabel metal2 s 121968 0 122024 400 6 s_axi_awaddr[10]
port 379 nsew signal output
rlabel metal2 s 126448 0 126504 400 6 s_axi_awaddr[11]
port 380 nsew signal output
rlabel metal2 s 130928 0 130984 400 6 s_axi_awaddr[12]
port 381 nsew signal output
rlabel metal2 s 135408 0 135464 400 6 s_axi_awaddr[13]
port 382 nsew signal output
rlabel metal2 s 139888 0 139944 400 6 s_axi_awaddr[14]
port 383 nsew signal output
rlabel metal2 s 144368 0 144424 400 6 s_axi_awaddr[15]
port 384 nsew signal output
rlabel metal2 s 148848 0 148904 400 6 s_axi_awaddr[16]
port 385 nsew signal output
rlabel metal2 s 153328 0 153384 400 6 s_axi_awaddr[17]
port 386 nsew signal output
rlabel metal2 s 157808 0 157864 400 6 s_axi_awaddr[18]
port 387 nsew signal output
rlabel metal2 s 162288 0 162344 400 6 s_axi_awaddr[19]
port 388 nsew signal output
rlabel metal2 s 53648 0 53704 400 6 s_axi_awaddr[1]
port 389 nsew signal output
rlabel metal2 s 166768 0 166824 400 6 s_axi_awaddr[20]
port 390 nsew signal output
rlabel metal2 s 171248 0 171304 400 6 s_axi_awaddr[21]
port 391 nsew signal output
rlabel metal2 s 175728 0 175784 400 6 s_axi_awaddr[22]
port 392 nsew signal output
rlabel metal2 s 180208 0 180264 400 6 s_axi_awaddr[23]
port 393 nsew signal output
rlabel metal2 s 184688 0 184744 400 6 s_axi_awaddr[24]
port 394 nsew signal output
rlabel metal2 s 189168 0 189224 400 6 s_axi_awaddr[25]
port 395 nsew signal output
rlabel metal2 s 193648 0 193704 400 6 s_axi_awaddr[26]
port 396 nsew signal output
rlabel metal2 s 198128 0 198184 400 6 s_axi_awaddr[27]
port 397 nsew signal output
rlabel metal2 s 202608 0 202664 400 6 s_axi_awaddr[28]
port 398 nsew signal output
rlabel metal2 s 207088 0 207144 400 6 s_axi_awaddr[29]
port 399 nsew signal output
rlabel metal2 s 67088 0 67144 400 6 s_axi_awaddr[2]
port 400 nsew signal output
rlabel metal2 s 211568 0 211624 400 6 s_axi_awaddr[30]
port 401 nsew signal output
rlabel metal2 s 216048 0 216104 400 6 s_axi_awaddr[31]
port 402 nsew signal output
rlabel metal2 s 78288 0 78344 400 6 s_axi_awaddr[3]
port 403 nsew signal output
rlabel metal2 s 87248 0 87304 400 6 s_axi_awaddr[4]
port 404 nsew signal output
rlabel metal2 s 93968 0 94024 400 6 s_axi_awaddr[5]
port 405 nsew signal output
rlabel metal2 s 100688 0 100744 400 6 s_axi_awaddr[6]
port 406 nsew signal output
rlabel metal2 s 107408 0 107464 400 6 s_axi_awaddr[7]
port 407 nsew signal output
rlabel metal2 s 113008 0 113064 400 6 s_axi_awaddr[8]
port 408 nsew signal output
rlabel metal2 s 117488 0 117544 400 6 s_axi_awaddr[9]
port 409 nsew signal output
rlabel metal2 s 40208 0 40264 400 6 s_axi_awburst[0]
port 410 nsew signal output
rlabel metal2 s 54768 0 54824 400 6 s_axi_awburst[1]
port 411 nsew signal output
rlabel metal2 s 41328 0 41384 400 6 s_axi_awcache[0]
port 412 nsew signal output
rlabel metal2 s 55888 0 55944 400 6 s_axi_awcache[1]
port 413 nsew signal output
rlabel metal2 s 68208 0 68264 400 6 s_axi_awcache[2]
port 414 nsew signal output
rlabel metal2 s 79408 0 79464 400 6 s_axi_awcache[3]
port 415 nsew signal output
rlabel metal2 s 17808 0 17864 400 6 s_axi_awid
port 416 nsew signal output
rlabel metal2 s 42448 0 42504 400 6 s_axi_awlen[0]
port 417 nsew signal output
rlabel metal2 s 57008 0 57064 400 6 s_axi_awlen[1]
port 418 nsew signal output
rlabel metal2 s 69328 0 69384 400 6 s_axi_awlen[2]
port 419 nsew signal output
rlabel metal2 s 80528 0 80584 400 6 s_axi_awlen[3]
port 420 nsew signal output
rlabel metal2 s 88368 0 88424 400 6 s_axi_awlen[4]
port 421 nsew signal output
rlabel metal2 s 95088 0 95144 400 6 s_axi_awlen[5]
port 422 nsew signal output
rlabel metal2 s 101808 0 101864 400 6 s_axi_awlen[6]
port 423 nsew signal output
rlabel metal2 s 108528 0 108584 400 6 s_axi_awlen[7]
port 424 nsew signal output
rlabel metal2 s 18928 0 18984 400 6 s_axi_awlock
port 425 nsew signal output
rlabel metal2 s 20048 0 20104 400 6 s_axi_awready
port 426 nsew signal input
rlabel metal2 s 43568 0 43624 400 6 s_axi_awsize[0]
port 427 nsew signal output
rlabel metal2 s 58128 0 58184 400 6 s_axi_awsize[1]
port 428 nsew signal output
rlabel metal2 s 70448 0 70504 400 6 s_axi_awsize[2]
port 429 nsew signal output
rlabel metal2 s 21168 0 21224 400 6 s_axi_awvalid
port 430 nsew signal output
rlabel metal2 s 22288 0 22344 400 6 s_axi_bid
port 431 nsew signal input
rlabel metal2 s 23408 0 23464 400 6 s_axi_bready
port 432 nsew signal output
rlabel metal2 s 24528 0 24584 400 6 s_axi_bvalid
port 433 nsew signal input
rlabel metal2 s 44688 0 44744 400 6 s_axi_rdata[0]
port 434 nsew signal input
rlabel metal2 s 123088 0 123144 400 6 s_axi_rdata[10]
port 435 nsew signal input
rlabel metal2 s 127568 0 127624 400 6 s_axi_rdata[11]
port 436 nsew signal input
rlabel metal2 s 132048 0 132104 400 6 s_axi_rdata[12]
port 437 nsew signal input
rlabel metal2 s 136528 0 136584 400 6 s_axi_rdata[13]
port 438 nsew signal input
rlabel metal2 s 141008 0 141064 400 6 s_axi_rdata[14]
port 439 nsew signal input
rlabel metal2 s 145488 0 145544 400 6 s_axi_rdata[15]
port 440 nsew signal input
rlabel metal2 s 149968 0 150024 400 6 s_axi_rdata[16]
port 441 nsew signal input
rlabel metal2 s 154448 0 154504 400 6 s_axi_rdata[17]
port 442 nsew signal input
rlabel metal2 s 158928 0 158984 400 6 s_axi_rdata[18]
port 443 nsew signal input
rlabel metal2 s 163408 0 163464 400 6 s_axi_rdata[19]
port 444 nsew signal input
rlabel metal2 s 59248 0 59304 400 6 s_axi_rdata[1]
port 445 nsew signal input
rlabel metal2 s 167888 0 167944 400 6 s_axi_rdata[20]
port 446 nsew signal input
rlabel metal2 s 172368 0 172424 400 6 s_axi_rdata[21]
port 447 nsew signal input
rlabel metal2 s 176848 0 176904 400 6 s_axi_rdata[22]
port 448 nsew signal input
rlabel metal2 s 181328 0 181384 400 6 s_axi_rdata[23]
port 449 nsew signal input
rlabel metal2 s 185808 0 185864 400 6 s_axi_rdata[24]
port 450 nsew signal input
rlabel metal2 s 190288 0 190344 400 6 s_axi_rdata[25]
port 451 nsew signal input
rlabel metal2 s 194768 0 194824 400 6 s_axi_rdata[26]
port 452 nsew signal input
rlabel metal2 s 199248 0 199304 400 6 s_axi_rdata[27]
port 453 nsew signal input
rlabel metal2 s 203728 0 203784 400 6 s_axi_rdata[28]
port 454 nsew signal input
rlabel metal2 s 208208 0 208264 400 6 s_axi_rdata[29]
port 455 nsew signal input
rlabel metal2 s 71568 0 71624 400 6 s_axi_rdata[2]
port 456 nsew signal input
rlabel metal2 s 212688 0 212744 400 6 s_axi_rdata[30]
port 457 nsew signal input
rlabel metal2 s 217168 0 217224 400 6 s_axi_rdata[31]
port 458 nsew signal input
rlabel metal2 s 81648 0 81704 400 6 s_axi_rdata[3]
port 459 nsew signal input
rlabel metal2 s 89488 0 89544 400 6 s_axi_rdata[4]
port 460 nsew signal input
rlabel metal2 s 96208 0 96264 400 6 s_axi_rdata[5]
port 461 nsew signal input
rlabel metal2 s 102928 0 102984 400 6 s_axi_rdata[6]
port 462 nsew signal input
rlabel metal2 s 109648 0 109704 400 6 s_axi_rdata[7]
port 463 nsew signal input
rlabel metal2 s 114128 0 114184 400 6 s_axi_rdata[8]
port 464 nsew signal input
rlabel metal2 s 118608 0 118664 400 6 s_axi_rdata[9]
port 465 nsew signal input
rlabel metal2 s 25648 0 25704 400 6 s_axi_rid
port 466 nsew signal input
rlabel metal2 s 26768 0 26824 400 6 s_axi_rlast
port 467 nsew signal input
rlabel metal2 s 27888 0 27944 400 6 s_axi_rready
port 468 nsew signal output
rlabel metal2 s 29008 0 29064 400 6 s_axi_rvalid
port 469 nsew signal input
rlabel metal2 s 45808 0 45864 400 6 s_axi_wdata[0]
port 470 nsew signal output
rlabel metal2 s 124208 0 124264 400 6 s_axi_wdata[10]
port 471 nsew signal output
rlabel metal2 s 128688 0 128744 400 6 s_axi_wdata[11]
port 472 nsew signal output
rlabel metal2 s 133168 0 133224 400 6 s_axi_wdata[12]
port 473 nsew signal output
rlabel metal2 s 137648 0 137704 400 6 s_axi_wdata[13]
port 474 nsew signal output
rlabel metal2 s 142128 0 142184 400 6 s_axi_wdata[14]
port 475 nsew signal output
rlabel metal2 s 146608 0 146664 400 6 s_axi_wdata[15]
port 476 nsew signal output
rlabel metal2 s 151088 0 151144 400 6 s_axi_wdata[16]
port 477 nsew signal output
rlabel metal2 s 155568 0 155624 400 6 s_axi_wdata[17]
port 478 nsew signal output
rlabel metal2 s 160048 0 160104 400 6 s_axi_wdata[18]
port 479 nsew signal output
rlabel metal2 s 164528 0 164584 400 6 s_axi_wdata[19]
port 480 nsew signal output
rlabel metal2 s 60368 0 60424 400 6 s_axi_wdata[1]
port 481 nsew signal output
rlabel metal2 s 169008 0 169064 400 6 s_axi_wdata[20]
port 482 nsew signal output
rlabel metal2 s 173488 0 173544 400 6 s_axi_wdata[21]
port 483 nsew signal output
rlabel metal2 s 177968 0 178024 400 6 s_axi_wdata[22]
port 484 nsew signal output
rlabel metal2 s 182448 0 182504 400 6 s_axi_wdata[23]
port 485 nsew signal output
rlabel metal2 s 186928 0 186984 400 6 s_axi_wdata[24]
port 486 nsew signal output
rlabel metal2 s 191408 0 191464 400 6 s_axi_wdata[25]
port 487 nsew signal output
rlabel metal2 s 195888 0 195944 400 6 s_axi_wdata[26]
port 488 nsew signal output
rlabel metal2 s 200368 0 200424 400 6 s_axi_wdata[27]
port 489 nsew signal output
rlabel metal2 s 204848 0 204904 400 6 s_axi_wdata[28]
port 490 nsew signal output
rlabel metal2 s 209328 0 209384 400 6 s_axi_wdata[29]
port 491 nsew signal output
rlabel metal2 s 72688 0 72744 400 6 s_axi_wdata[2]
port 492 nsew signal output
rlabel metal2 s 213808 0 213864 400 6 s_axi_wdata[30]
port 493 nsew signal output
rlabel metal2 s 218288 0 218344 400 6 s_axi_wdata[31]
port 494 nsew signal output
rlabel metal2 s 82768 0 82824 400 6 s_axi_wdata[3]
port 495 nsew signal output
rlabel metal2 s 90608 0 90664 400 6 s_axi_wdata[4]
port 496 nsew signal output
rlabel metal2 s 97328 0 97384 400 6 s_axi_wdata[5]
port 497 nsew signal output
rlabel metal2 s 104048 0 104104 400 6 s_axi_wdata[6]
port 498 nsew signal output
rlabel metal2 s 110768 0 110824 400 6 s_axi_wdata[7]
port 499 nsew signal output
rlabel metal2 s 115248 0 115304 400 6 s_axi_wdata[8]
port 500 nsew signal output
rlabel metal2 s 119728 0 119784 400 6 s_axi_wdata[9]
port 501 nsew signal output
rlabel metal2 s 30128 0 30184 400 6 s_axi_wlast
port 502 nsew signal output
rlabel metal2 s 31248 0 31304 400 6 s_axi_wready
port 503 nsew signal input
rlabel metal2 s 46928 0 46984 400 6 s_axi_wstrb[0]
port 504 nsew signal output
rlabel metal2 s 61488 0 61544 400 6 s_axi_wstrb[1]
port 505 nsew signal output
rlabel metal2 s 73808 0 73864 400 6 s_axi_wstrb[2]
port 506 nsew signal output
rlabel metal2 s 83888 0 83944 400 6 s_axi_wstrb[3]
port 507 nsew signal output
rlabel metal2 s 32368 0 32424 400 6 s_axi_wvalid
port 508 nsew signal output
rlabel metal4 s 2224 1538 2384 298342 6 vdd
port 509 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 298342 6 vdd
port 509 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 298342 6 vdd
port 509 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 298342 6 vdd
port 509 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 298342 6 vdd
port 509 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 298342 6 vdd
port 509 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 298342 6 vdd
port 509 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 298342 6 vdd
port 509 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 298342 6 vdd
port 509 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 298342 6 vdd
port 509 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 298342 6 vdd
port 509 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 298342 6 vdd
port 509 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 298342 6 vdd
port 509 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 298342 6 vdd
port 509 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 298342 6 vdd
port 509 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 298342 6 vdd
port 509 nsew power bidirectional
rlabel metal4 s 247984 1538 248144 298342 6 vdd
port 509 nsew power bidirectional
rlabel metal4 s 263344 1538 263504 298342 6 vdd
port 509 nsew power bidirectional
rlabel metal4 s 278704 1538 278864 298342 6 vdd
port 509 nsew power bidirectional
rlabel metal4 s 294064 1538 294224 298342 6 vdd
port 509 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 298342 6 vss
port 510 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 298342 6 vss
port 510 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 298342 6 vss
port 510 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 298342 6 vss
port 510 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 298342 6 vss
port 510 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 298342 6 vss
port 510 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 298342 6 vss
port 510 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 298342 6 vss
port 510 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 298342 6 vss
port 510 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 298342 6 vss
port 510 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 298342 6 vss
port 510 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 298342 6 vss
port 510 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 298342 6 vss
port 510 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 298342 6 vss
port 510 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 298342 6 vss
port 510 nsew ground bidirectional
rlabel metal4 s 240304 1538 240464 298342 6 vss
port 510 nsew ground bidirectional
rlabel metal4 s 255664 1538 255824 298342 6 vss
port 510 nsew ground bidirectional
rlabel metal4 s 271024 1538 271184 298342 6 vss
port 510 nsew ground bidirectional
rlabel metal4 s 286384 1538 286544 298342 6 vss
port 510 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 300000 300000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 356298322
string GDS_FILE /home/m/Builds/caravel_user_project/openlane/SoC/runs/23_11_30_13_33/results/signoff/SoC.magic.gds
string GDS_START 208484
<< end >>

