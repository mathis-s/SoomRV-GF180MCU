VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO SoC
  CLASS BLOCK ;
  FOREIGN SoC ;
  ORIGIN 0.000 0.000 ;
  SIZE 3000.000 BY 3000.000 ;
  PIN IN_DCT_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.399000 ;
    ANTENNADIFFAREA 1.641600 ;
    PORT
      LAYER Metal2 ;
        RECT 469.280 2996.000 469.840 3000.000 ;
    END
  END IN_DCT_data[0]
  PIN IN_DCT_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.096500 ;
    ANTENNADIFFAREA 1.231200 ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 2996.000 245.840 3000.000 ;
    END
  END IN_DCT_data[10]
  PIN IN_DCT_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.692000 ;
    ANTENNADIFFAREA 1.641600 ;
    PORT
      LAYER Metal2 ;
        RECT 222.880 2996.000 223.440 3000.000 ;
    END
  END IN_DCT_data[11]
  PIN IN_DCT_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.694500 ;
    ANTENNADIFFAREA 1.641600 ;
    PORT
      LAYER Metal2 ;
        RECT 200.480 2996.000 201.040 3000.000 ;
    END
  END IN_DCT_data[12]
  PIN IN_DCT_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.445000 ;
    ANTENNADIFFAREA 1.231200 ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 2996.000 178.640 3000.000 ;
    END
  END IN_DCT_data[13]
  PIN IN_DCT_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.955500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 2996.000 156.240 3000.000 ;
    END
  END IN_DCT_data[14]
  PIN IN_DCT_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.643500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 133.280 2996.000 133.840 3000.000 ;
    END
  END IN_DCT_data[15]
  PIN IN_DCT_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.794000 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 2996.000 111.440 3000.000 ;
    END
  END IN_DCT_data[16]
  PIN IN_DCT_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.694500 ;
    ANTENNADIFFAREA 1.641600 ;
    PORT
      LAYER Metal2 ;
        RECT 88.480 2996.000 89.040 3000.000 ;
    END
  END IN_DCT_data[17]
  PIN IN_DCT_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.598000 ;
    ANTENNADIFFAREA 1.231200 ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 2996.000 66.640 3000.000 ;
    END
  END IN_DCT_data[18]
  PIN IN_DCT_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.694500 ;
    ANTENNADIFFAREA 1.641600 ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 2996.000 44.240 3000.000 ;
    END
  END IN_DCT_data[19]
  PIN IN_DCT_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.796500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 446.880 2996.000 447.440 3000.000 ;
    END
  END IN_DCT_data[1]
  PIN IN_DCT_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.697500 ;
    ANTENNADIFFAREA 1.641600 ;
    PORT
      LAYER Metal2 ;
        RECT 21.280 2996.000 21.840 3000.000 ;
    END
  END IN_DCT_data[20]
  PIN IN_DCT_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.796500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 424.480 2996.000 425.040 3000.000 ;
    END
  END IN_DCT_data[2]
  PIN IN_DCT_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000500 ;
    ANTENNADIFFAREA 1.641600 ;
    PORT
      LAYER Metal2 ;
        RECT 402.080 2996.000 402.640 3000.000 ;
    END
  END IN_DCT_data[3]
  PIN IN_DCT_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.196000 ;
    ANTENNADIFFAREA 1.641600 ;
    PORT
      LAYER Metal2 ;
        RECT 379.680 2996.000 380.240 3000.000 ;
    END
  END IN_DCT_data[4]
  PIN IN_DCT_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.592500 ;
    ANTENNADIFFAREA 1.231200 ;
    PORT
      LAYER Metal2 ;
        RECT 357.280 2996.000 357.840 3000.000 ;
    END
  END IN_DCT_data[5]
  PIN IN_DCT_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.553000 ;
    ANTENNADIFFAREA 1.231200 ;
    PORT
      LAYER Metal2 ;
        RECT 334.880 2996.000 335.440 3000.000 ;
    END
  END IN_DCT_data[6]
  PIN IN_DCT_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.595500 ;
    ANTENNADIFFAREA 1.231200 ;
    PORT
      LAYER Metal2 ;
        RECT 312.480 2996.000 313.040 3000.000 ;
    END
  END IN_DCT_data[7]
  PIN IN_DCT_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.700000 ;
    ANTENNADIFFAREA 1.641600 ;
    PORT
      LAYER Metal2 ;
        RECT 290.080 2996.000 290.640 3000.000 ;
    END
  END IN_DCT_data[8]
  PIN IN_DCT_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.000000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 267.680 2996.000 268.240 3000.000 ;
    END
  END IN_DCT_data[9]
  PIN IN_DC_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1902.880 2996.000 1903.440 3000.000 ;
    END
  END IN_DC_data[0]
  PIN IN_DC_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1678.880 2996.000 1679.440 3000.000 ;
    END
  END IN_DC_data[10]
  PIN IN_DC_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 1656.480 2996.000 1657.040 3000.000 ;
    END
  END IN_DC_data[11]
  PIN IN_DC_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1634.080 2996.000 1634.640 3000.000 ;
    END
  END IN_DC_data[12]
  PIN IN_DC_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1611.680 2996.000 1612.240 3000.000 ;
    END
  END IN_DC_data[13]
  PIN IN_DC_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1589.280 2996.000 1589.840 3000.000 ;
    END
  END IN_DC_data[14]
  PIN IN_DC_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1566.880 2996.000 1567.440 3000.000 ;
    END
  END IN_DC_data[15]
  PIN IN_DC_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 1544.480 2996.000 1545.040 3000.000 ;
    END
  END IN_DC_data[16]
  PIN IN_DC_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1522.080 2996.000 1522.640 3000.000 ;
    END
  END IN_DC_data[17]
  PIN IN_DC_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1499.680 2996.000 1500.240 3000.000 ;
    END
  END IN_DC_data[18]
  PIN IN_DC_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1477.280 2996.000 1477.840 3000.000 ;
    END
  END IN_DC_data[19]
  PIN IN_DC_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1880.480 2996.000 1881.040 3000.000 ;
    END
  END IN_DC_data[1]
  PIN IN_DC_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1454.880 2996.000 1455.440 3000.000 ;
    END
  END IN_DC_data[20]
  PIN IN_DC_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1432.480 2996.000 1433.040 3000.000 ;
    END
  END IN_DC_data[21]
  PIN IN_DC_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1410.080 2996.000 1410.640 3000.000 ;
    END
  END IN_DC_data[22]
  PIN IN_DC_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1387.680 2996.000 1388.240 3000.000 ;
    END
  END IN_DC_data[23]
  PIN IN_DC_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 1365.280 2996.000 1365.840 3000.000 ;
    END
  END IN_DC_data[24]
  PIN IN_DC_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1342.880 2996.000 1343.440 3000.000 ;
    END
  END IN_DC_data[25]
  PIN IN_DC_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1320.480 2996.000 1321.040 3000.000 ;
    END
  END IN_DC_data[26]
  PIN IN_DC_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1298.080 2996.000 1298.640 3000.000 ;
    END
  END IN_DC_data[27]
  PIN IN_DC_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1275.680 2996.000 1276.240 3000.000 ;
    END
  END IN_DC_data[28]
  PIN IN_DC_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1253.280 2996.000 1253.840 3000.000 ;
    END
  END IN_DC_data[29]
  PIN IN_DC_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1858.080 2996.000 1858.640 3000.000 ;
    END
  END IN_DC_data[2]
  PIN IN_DC_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1230.880 2996.000 1231.440 3000.000 ;
    END
  END IN_DC_data[30]
  PIN IN_DC_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1208.480 2996.000 1209.040 3000.000 ;
    END
  END IN_DC_data[31]
  PIN IN_DC_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1835.680 2996.000 1836.240 3000.000 ;
    END
  END IN_DC_data[3]
  PIN IN_DC_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1813.280 2996.000 1813.840 3000.000 ;
    END
  END IN_DC_data[4]
  PIN IN_DC_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1790.880 2996.000 1791.440 3000.000 ;
    END
  END IN_DC_data[5]
  PIN IN_DC_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1768.480 2996.000 1769.040 3000.000 ;
    END
  END IN_DC_data[6]
  PIN IN_DC_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1746.080 2996.000 1746.640 3000.000 ;
    END
  END IN_DC_data[7]
  PIN IN_DC_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1723.680 2996.000 1724.240 3000.000 ;
    END
  END IN_DC_data[8]
  PIN IN_DC_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1701.280 2996.000 1701.840 3000.000 ;
    END
  END IN_DC_data[9]
  PIN IN_ICT_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 502.880 4.000 503.440 ;
    END
  END IN_ICT_data[0]
  PIN IN_ICT_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.159000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 278.880 4.000 279.440 ;
    END
  END IN_ICT_data[10]
  PIN IN_ICT_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.598000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 256.480 4.000 257.040 ;
    END
  END IN_ICT_data[11]
  PIN IN_ICT_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.135500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 234.080 4.000 234.640 ;
    END
  END IN_ICT_data[12]
  PIN IN_ICT_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.006000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 211.680 4.000 212.240 ;
    END
  END IN_ICT_data[13]
  PIN IN_ICT_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.598000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 189.280 4.000 189.840 ;
    END
  END IN_ICT_data[14]
  PIN IN_ICT_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.598000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 166.880 4.000 167.440 ;
    END
  END IN_ICT_data[15]
  PIN IN_ICT_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.159000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 144.480 4.000 145.040 ;
    END
  END IN_ICT_data[16]
  PIN IN_ICT_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.198500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 122.080 4.000 122.640 ;
    END
  END IN_ICT_data[17]
  PIN IN_ICT_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.159000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 99.680 4.000 100.240 ;
    END
  END IN_ICT_data[18]
  PIN IN_ICT_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.201500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 77.280 4.000 77.840 ;
    END
  END IN_ICT_data[19]
  PIN IN_ICT_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.198500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 480.480 4.000 481.040 ;
    END
  END IN_ICT_data[1]
  PIN IN_ICT_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.198500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 54.880 4.000 55.440 ;
    END
  END IN_ICT_data[20]
  PIN IN_ICT_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.198500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 458.080 4.000 458.640 ;
    END
  END IN_ICT_data[2]
  PIN IN_ICT_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.598000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 435.680 4.000 436.240 ;
    END
  END IN_ICT_data[3]
  PIN IN_ICT_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.201500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 413.280 4.000 413.840 ;
    END
  END IN_ICT_data[4]
  PIN IN_ICT_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.982500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 390.880 4.000 391.440 ;
    END
  END IN_ICT_data[5]
  PIN IN_ICT_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.198500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 368.480 4.000 369.040 ;
    END
  END IN_ICT_data[6]
  PIN IN_ICT_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.159000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 346.080 4.000 346.640 ;
    END
  END IN_ICT_data[7]
  PIN IN_ICT_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.159000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 323.680 4.000 324.240 ;
    END
  END IN_ICT_data[8]
  PIN IN_ICT_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.198500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 301.280 4.000 301.840 ;
    END
  END IN_ICT_data[9]
  PIN IN_IC_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1936.480 4.000 1937.040 ;
    END
  END IN_IC_data[0]
  PIN IN_IC_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1712.480 4.000 1713.040 ;
    END
  END IN_IC_data[10]
  PIN IN_IC_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1690.080 4.000 1690.640 ;
    END
  END IN_IC_data[11]
  PIN IN_IC_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1667.680 4.000 1668.240 ;
    END
  END IN_IC_data[12]
  PIN IN_IC_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1645.280 4.000 1645.840 ;
    END
  END IN_IC_data[13]
  PIN IN_IC_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1622.880 4.000 1623.440 ;
    END
  END IN_IC_data[14]
  PIN IN_IC_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1600.480 4.000 1601.040 ;
    END
  END IN_IC_data[15]
  PIN IN_IC_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1578.080 4.000 1578.640 ;
    END
  END IN_IC_data[16]
  PIN IN_IC_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1555.680 4.000 1556.240 ;
    END
  END IN_IC_data[17]
  PIN IN_IC_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1533.280 4.000 1533.840 ;
    END
  END IN_IC_data[18]
  PIN IN_IC_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1510.880 4.000 1511.440 ;
    END
  END IN_IC_data[19]
  PIN IN_IC_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1914.080 4.000 1914.640 ;
    END
  END IN_IC_data[1]
  PIN IN_IC_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1488.480 4.000 1489.040 ;
    END
  END IN_IC_data[20]
  PIN IN_IC_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1466.080 4.000 1466.640 ;
    END
  END IN_IC_data[21]
  PIN IN_IC_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1443.680 4.000 1444.240 ;
    END
  END IN_IC_data[22]
  PIN IN_IC_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1421.280 4.000 1421.840 ;
    END
  END IN_IC_data[23]
  PIN IN_IC_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1398.880 4.000 1399.440 ;
    END
  END IN_IC_data[24]
  PIN IN_IC_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1376.480 4.000 1377.040 ;
    END
  END IN_IC_data[25]
  PIN IN_IC_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1354.080 4.000 1354.640 ;
    END
  END IN_IC_data[26]
  PIN IN_IC_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1331.680 4.000 1332.240 ;
    END
  END IN_IC_data[27]
  PIN IN_IC_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1309.280 4.000 1309.840 ;
    END
  END IN_IC_data[28]
  PIN IN_IC_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1286.880 4.000 1287.440 ;
    END
  END IN_IC_data[29]
  PIN IN_IC_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1891.680 4.000 1892.240 ;
    END
  END IN_IC_data[2]
  PIN IN_IC_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1264.480 4.000 1265.040 ;
    END
  END IN_IC_data[30]
  PIN IN_IC_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1242.080 4.000 1242.640 ;
    END
  END IN_IC_data[31]
  PIN IN_IC_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1869.280 4.000 1869.840 ;
    END
  END IN_IC_data[3]
  PIN IN_IC_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1846.880 4.000 1847.440 ;
    END
  END IN_IC_data[4]
  PIN IN_IC_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1824.480 4.000 1825.040 ;
    END
  END IN_IC_data[5]
  PIN IN_IC_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1802.080 4.000 1802.640 ;
    END
  END IN_IC_data[6]
  PIN IN_IC_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1779.680 4.000 1780.240 ;
    END
  END IN_IC_data[7]
  PIN IN_IC_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1757.280 4.000 1757.840 ;
    END
  END IN_IC_data[8]
  PIN IN_IC_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1734.880 4.000 1735.440 ;
    END
  END IN_IC_data[9]
  PIN OUT_DCT_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.055600 ;
    PORT
      LAYER Metal2 ;
        RECT 1118.880 2996.000 1119.440 3000.000 ;
    END
  END OUT_DCT_addr[0]
  PIN OUT_DCT_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.055600 ;
    PORT
      LAYER Metal2 ;
        RECT 1074.080 2996.000 1074.640 3000.000 ;
    END
  END OUT_DCT_addr[1]
  PIN OUT_DCT_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.055600 ;
    PORT
      LAYER Metal2 ;
        RECT 1029.280 2996.000 1029.840 3000.000 ;
    END
  END OUT_DCT_addr[2]
  PIN OUT_DCT_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.055600 ;
    PORT
      LAYER Metal2 ;
        RECT 984.480 2996.000 985.040 3000.000 ;
    END
  END OUT_DCT_addr[3]
  PIN OUT_DCT_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.055600 ;
    PORT
      LAYER Metal2 ;
        RECT 939.680 2996.000 940.240 3000.000 ;
    END
  END OUT_DCT_addr[4]
  PIN OUT_DCT_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.948400 ;
    PORT
      LAYER Metal2 ;
        RECT 894.880 2996.000 895.440 3000.000 ;
    END
  END OUT_DCT_addr[5]
  PIN OUT_DCT_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.055600 ;
    PORT
      LAYER Metal2 ;
        RECT 850.080 2996.000 850.640 3000.000 ;
    END
  END OUT_DCT_addr[6]
  PIN OUT_DCT_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.055600 ;
    PORT
      LAYER Metal2 ;
        RECT 805.280 2996.000 805.840 3000.000 ;
    END
  END OUT_DCT_addr[7]
  PIN OUT_DCT_ce
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1186.080 2996.000 1186.640 3000.000 ;
    END
  END OUT_DCT_ce
  PIN OUT_DCT_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1096.480 2996.000 1097.040 3000.000 ;
    END
  END OUT_DCT_data[0]
  PIN OUT_DCT_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal2 ;
        RECT 715.680 2996.000 716.240 3000.000 ;
    END
  END OUT_DCT_data[10]
  PIN OUT_DCT_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal2 ;
        RECT 693.280 2996.000 693.840 3000.000 ;
    END
  END OUT_DCT_data[11]
  PIN OUT_DCT_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal2 ;
        RECT 670.880 2996.000 671.440 3000.000 ;
    END
  END OUT_DCT_data[12]
  PIN OUT_DCT_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal2 ;
        RECT 648.480 2996.000 649.040 3000.000 ;
    END
  END OUT_DCT_data[13]
  PIN OUT_DCT_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal2 ;
        RECT 626.080 2996.000 626.640 3000.000 ;
    END
  END OUT_DCT_data[14]
  PIN OUT_DCT_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal2 ;
        RECT 603.680 2996.000 604.240 3000.000 ;
    END
  END OUT_DCT_data[15]
  PIN OUT_DCT_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal2 ;
        RECT 581.280 2996.000 581.840 3000.000 ;
    END
  END OUT_DCT_data[16]
  PIN OUT_DCT_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal2 ;
        RECT 558.880 2996.000 559.440 3000.000 ;
    END
  END OUT_DCT_data[17]
  PIN OUT_DCT_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal2 ;
        RECT 536.480 2996.000 537.040 3000.000 ;
    END
  END OUT_DCT_data[18]
  PIN OUT_DCT_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal2 ;
        RECT 514.080 2996.000 514.640 3000.000 ;
    END
  END OUT_DCT_data[19]
  PIN OUT_DCT_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal2 ;
        RECT 1051.680 2996.000 1052.240 3000.000 ;
    END
  END OUT_DCT_data[1]
  PIN OUT_DCT_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal2 ;
        RECT 491.680 2996.000 492.240 3000.000 ;
    END
  END OUT_DCT_data[20]
  PIN OUT_DCT_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal2 ;
        RECT 1006.880 2996.000 1007.440 3000.000 ;
    END
  END OUT_DCT_data[2]
  PIN OUT_DCT_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal2 ;
        RECT 962.080 2996.000 962.640 3000.000 ;
    END
  END OUT_DCT_data[3]
  PIN OUT_DCT_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal2 ;
        RECT 917.280 2996.000 917.840 3000.000 ;
    END
  END OUT_DCT_data[4]
  PIN OUT_DCT_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal2 ;
        RECT 872.480 2996.000 873.040 3000.000 ;
    END
  END OUT_DCT_data[5]
  PIN OUT_DCT_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal2 ;
        RECT 827.680 2996.000 828.240 3000.000 ;
    END
  END OUT_DCT_data[6]
  PIN OUT_DCT_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal2 ;
        RECT 782.880 2996.000 783.440 3000.000 ;
    END
  END OUT_DCT_data[7]
  PIN OUT_DCT_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal2 ;
        RECT 760.480 2996.000 761.040 3000.000 ;
    END
  END OUT_DCT_data[8]
  PIN OUT_DCT_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal2 ;
        RECT 738.080 2996.000 738.640 3000.000 ;
    END
  END OUT_DCT_data[9]
  PIN OUT_DCT_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.593500 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1163.680 2996.000 1164.240 3000.000 ;
    END
  END OUT_DCT_we
  PIN OUT_DCT_wm
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1141.280 2996.000 1141.840 3000.000 ;
    END
  END OUT_DCT_wm
  PIN OUT_DC_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 2933.280 2996.000 2933.840 3000.000 ;
    END
  END OUT_DC_addr[0]
  PIN OUT_DC_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 2866.080 2996.000 2866.640 3000.000 ;
    END
  END OUT_DC_addr[1]
  PIN OUT_DC_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2798.880 2996.000 2799.440 3000.000 ;
    END
  END OUT_DC_addr[2]
  PIN OUT_DC_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2731.680 2996.000 2732.240 3000.000 ;
    END
  END OUT_DC_addr[3]
  PIN OUT_DC_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2664.480 2996.000 2665.040 3000.000 ;
    END
  END OUT_DC_addr[4]
  PIN OUT_DC_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2619.680 2996.000 2620.240 3000.000 ;
    END
  END OUT_DC_addr[5]
  PIN OUT_DC_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2574.880 2996.000 2575.440 3000.000 ;
    END
  END OUT_DC_addr[6]
  PIN OUT_DC_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2530.080 2996.000 2530.640 3000.000 ;
    END
  END OUT_DC_addr[7]
  PIN OUT_DC_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2485.280 2996.000 2485.840 3000.000 ;
    END
  END OUT_DC_addr[8]
  PIN OUT_DC_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.145600 ;
    PORT
      LAYER Metal2 ;
        RECT 2440.480 2996.000 2441.040 3000.000 ;
    END
  END OUT_DC_addr[9]
  PIN OUT_DC_ce
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2978.080 2996.000 2978.640 3000.000 ;
    END
  END OUT_DC_ce
  PIN OUT_DC_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.259900 ;
    PORT
      LAYER Metal2 ;
        RECT 2910.880 2996.000 2911.440 3000.000 ;
    END
  END OUT_DC_data[0]
  PIN OUT_DC_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2395.680 2996.000 2396.240 3000.000 ;
    END
  END OUT_DC_data[10]
  PIN OUT_DC_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2373.280 2996.000 2373.840 3000.000 ;
    END
  END OUT_DC_data[11]
  PIN OUT_DC_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2350.880 2996.000 2351.440 3000.000 ;
    END
  END OUT_DC_data[12]
  PIN OUT_DC_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2328.480 2996.000 2329.040 3000.000 ;
    END
  END OUT_DC_data[13]
  PIN OUT_DC_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2306.080 2996.000 2306.640 3000.000 ;
    END
  END OUT_DC_data[14]
  PIN OUT_DC_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2283.680 2996.000 2284.240 3000.000 ;
    END
  END OUT_DC_data[15]
  PIN OUT_DC_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2261.280 2996.000 2261.840 3000.000 ;
    END
  END OUT_DC_data[16]
  PIN OUT_DC_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2238.880 2996.000 2239.440 3000.000 ;
    END
  END OUT_DC_data[17]
  PIN OUT_DC_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2216.480 2996.000 2217.040 3000.000 ;
    END
  END OUT_DC_data[18]
  PIN OUT_DC_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2194.080 2996.000 2194.640 3000.000 ;
    END
  END OUT_DC_data[19]
  PIN OUT_DC_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.259900 ;
    PORT
      LAYER Metal2 ;
        RECT 2843.680 2996.000 2844.240 3000.000 ;
    END
  END OUT_DC_data[1]
  PIN OUT_DC_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2171.680 2996.000 2172.240 3000.000 ;
    END
  END OUT_DC_data[20]
  PIN OUT_DC_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2149.280 2996.000 2149.840 3000.000 ;
    END
  END OUT_DC_data[21]
  PIN OUT_DC_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2126.880 2996.000 2127.440 3000.000 ;
    END
  END OUT_DC_data[22]
  PIN OUT_DC_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2104.480 2996.000 2105.040 3000.000 ;
    END
  END OUT_DC_data[23]
  PIN OUT_DC_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2082.080 2996.000 2082.640 3000.000 ;
    END
  END OUT_DC_data[24]
  PIN OUT_DC_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2059.680 2996.000 2060.240 3000.000 ;
    END
  END OUT_DC_data[25]
  PIN OUT_DC_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2037.280 2996.000 2037.840 3000.000 ;
    END
  END OUT_DC_data[26]
  PIN OUT_DC_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2014.880 2996.000 2015.440 3000.000 ;
    END
  END OUT_DC_data[27]
  PIN OUT_DC_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1992.480 2996.000 1993.040 3000.000 ;
    END
  END OUT_DC_data[28]
  PIN OUT_DC_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1970.080 2996.000 1970.640 3000.000 ;
    END
  END OUT_DC_data[29]
  PIN OUT_DC_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.259900 ;
    PORT
      LAYER Metal2 ;
        RECT 2776.480 2996.000 2777.040 3000.000 ;
    END
  END OUT_DC_data[2]
  PIN OUT_DC_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1947.680 2996.000 1948.240 3000.000 ;
    END
  END OUT_DC_data[30]
  PIN OUT_DC_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1925.280 2996.000 1925.840 3000.000 ;
    END
  END OUT_DC_data[31]
  PIN OUT_DC_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.259900 ;
    PORT
      LAYER Metal2 ;
        RECT 2709.280 2996.000 2709.840 3000.000 ;
    END
  END OUT_DC_data[3]
  PIN OUT_DC_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.259900 ;
    PORT
      LAYER Metal2 ;
        RECT 2642.080 2996.000 2642.640 3000.000 ;
    END
  END OUT_DC_data[4]
  PIN OUT_DC_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.259900 ;
    PORT
      LAYER Metal2 ;
        RECT 2597.280 2996.000 2597.840 3000.000 ;
    END
  END OUT_DC_data[5]
  PIN OUT_DC_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.259900 ;
    PORT
      LAYER Metal2 ;
        RECT 2552.480 2996.000 2553.040 3000.000 ;
    END
  END OUT_DC_data[6]
  PIN OUT_DC_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.259900 ;
    PORT
      LAYER Metal2 ;
        RECT 2507.680 2996.000 2508.240 3000.000 ;
    END
  END OUT_DC_data[7]
  PIN OUT_DC_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.259900 ;
    PORT
      LAYER Metal2 ;
        RECT 2462.880 2996.000 2463.440 3000.000 ;
    END
  END OUT_DC_data[8]
  PIN OUT_DC_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2418.080 2996.000 2418.640 3000.000 ;
    END
  END OUT_DC_data[9]
  PIN OUT_DC_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.291500 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2955.680 2996.000 2956.240 3000.000 ;
    END
  END OUT_DC_we
  PIN OUT_DC_wm[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal2 ;
        RECT 2888.480 2996.000 2889.040 3000.000 ;
    END
  END OUT_DC_wm[0]
  PIN OUT_DC_wm[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal2 ;
        RECT 2821.280 2996.000 2821.840 3000.000 ;
    END
  END OUT_DC_wm[1]
  PIN OUT_DC_wm[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal2 ;
        RECT 2754.080 2996.000 2754.640 3000.000 ;
    END
  END OUT_DC_wm[2]
  PIN OUT_DC_wm[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal2 ;
        RECT 2686.880 2996.000 2687.440 3000.000 ;
    END
  END OUT_DC_wm[3]
  PIN OUT_ICT_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.489200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1152.480 4.000 1153.040 ;
    END
  END OUT_ICT_addr[0]
  PIN OUT_ICT_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.145600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1107.680 4.000 1108.240 ;
    END
  END OUT_ICT_addr[1]
  PIN OUT_ICT_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.145600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1062.880 4.000 1063.440 ;
    END
  END OUT_ICT_addr[2]
  PIN OUT_ICT_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.145600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1018.080 4.000 1018.640 ;
    END
  END OUT_ICT_addr[3]
  PIN OUT_ICT_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.988400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 973.280 4.000 973.840 ;
    END
  END OUT_ICT_addr[4]
  PIN OUT_ICT_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.145600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 928.480 4.000 929.040 ;
    END
  END OUT_ICT_addr[5]
  PIN OUT_ICT_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.988400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 883.680 4.000 884.240 ;
    END
  END OUT_ICT_addr[6]
  PIN OUT_ICT_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.145600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 838.880 4.000 839.440 ;
    END
  END OUT_ICT_addr[7]
  PIN OUT_ICT_ce
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.983200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1219.680 4.000 1220.240 ;
    END
  END OUT_ICT_ce
  PIN OUT_ICT_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.914000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1130.080 4.000 1130.640 ;
    END
  END OUT_ICT_data[0]
  PIN OUT_ICT_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 749.280 4.000 749.840 ;
    END
  END OUT_ICT_data[10]
  PIN OUT_ICT_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 726.880 4.000 727.440 ;
    END
  END OUT_ICT_data[11]
  PIN OUT_ICT_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 704.480 4.000 705.040 ;
    END
  END OUT_ICT_data[12]
  PIN OUT_ICT_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 682.080 4.000 682.640 ;
    END
  END OUT_ICT_data[13]
  PIN OUT_ICT_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 659.680 4.000 660.240 ;
    END
  END OUT_ICT_data[14]
  PIN OUT_ICT_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 637.280 4.000 637.840 ;
    END
  END OUT_ICT_data[15]
  PIN OUT_ICT_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 614.880 4.000 615.440 ;
    END
  END OUT_ICT_data[16]
  PIN OUT_ICT_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 592.480 4.000 593.040 ;
    END
  END OUT_ICT_data[17]
  PIN OUT_ICT_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 570.080 4.000 570.640 ;
    END
  END OUT_ICT_data[18]
  PIN OUT_ICT_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 547.680 4.000 548.240 ;
    END
  END OUT_ICT_data[19]
  PIN OUT_ICT_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1085.280 4.000 1085.840 ;
    END
  END OUT_ICT_data[1]
  PIN OUT_ICT_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 525.280 4.000 525.840 ;
    END
  END OUT_ICT_data[20]
  PIN OUT_ICT_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1040.480 4.000 1041.040 ;
    END
  END OUT_ICT_data[2]
  PIN OUT_ICT_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 995.680 4.000 996.240 ;
    END
  END OUT_ICT_data[3]
  PIN OUT_ICT_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 950.880 4.000 951.440 ;
    END
  END OUT_ICT_data[4]
  PIN OUT_ICT_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 906.080 4.000 906.640 ;
    END
  END OUT_ICT_data[5]
  PIN OUT_ICT_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 861.280 4.000 861.840 ;
    END
  END OUT_ICT_data[6]
  PIN OUT_ICT_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 816.480 4.000 817.040 ;
    END
  END OUT_ICT_data[7]
  PIN OUT_ICT_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 794.080 4.000 794.640 ;
    END
  END OUT_ICT_data[8]
  PIN OUT_ICT_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 771.680 4.000 772.240 ;
    END
  END OUT_ICT_data[9]
  PIN OUT_ICT_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.497500 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1197.280 4.000 1197.840 ;
    END
  END OUT_ICT_we
  PIN OUT_ICT_wm
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1174.880 4.000 1175.440 ;
    END
  END OUT_ICT_wm
  PIN OUT_IC_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2877.280 4.000 2877.840 ;
    END
  END OUT_IC_addr[0]
  PIN OUT_IC_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2832.480 4.000 2833.040 ;
    END
  END OUT_IC_addr[1]
  PIN OUT_IC_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2787.680 4.000 2788.240 ;
    END
  END OUT_IC_addr[2]
  PIN OUT_IC_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2742.880 4.000 2743.440 ;
    END
  END OUT_IC_addr[3]
  PIN OUT_IC_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2698.080 4.000 2698.640 ;
    END
  END OUT_IC_addr[4]
  PIN OUT_IC_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.988400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2653.280 4.000 2653.840 ;
    END
  END OUT_IC_addr[5]
  PIN OUT_IC_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.988400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2608.480 4.000 2609.040 ;
    END
  END OUT_IC_addr[6]
  PIN OUT_IC_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2563.680 4.000 2564.240 ;
    END
  END OUT_IC_addr[7]
  PIN OUT_IC_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2518.880 4.000 2519.440 ;
    END
  END OUT_IC_addr[8]
  PIN OUT_IC_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2474.080 4.000 2474.640 ;
    END
  END OUT_IC_addr[9]
  PIN OUT_IC_ce
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2944.480 4.000 2945.040 ;
    END
  END OUT_IC_ce
  PIN OUT_IC_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2854.880 4.000 2855.440 ;
    END
  END OUT_IC_data[0]
  PIN OUT_IC_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2429.280 4.000 2429.840 ;
    END
  END OUT_IC_data[10]
  PIN OUT_IC_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2406.880 4.000 2407.440 ;
    END
  END OUT_IC_data[11]
  PIN OUT_IC_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2384.480 4.000 2385.040 ;
    END
  END OUT_IC_data[12]
  PIN OUT_IC_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2362.080 4.000 2362.640 ;
    END
  END OUT_IC_data[13]
  PIN OUT_IC_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2339.680 4.000 2340.240 ;
    END
  END OUT_IC_data[14]
  PIN OUT_IC_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2317.280 4.000 2317.840 ;
    END
  END OUT_IC_data[15]
  PIN OUT_IC_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2294.880 4.000 2295.440 ;
    END
  END OUT_IC_data[16]
  PIN OUT_IC_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2272.480 4.000 2273.040 ;
    END
  END OUT_IC_data[17]
  PIN OUT_IC_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2250.080 4.000 2250.640 ;
    END
  END OUT_IC_data[18]
  PIN OUT_IC_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2227.680 4.000 2228.240 ;
    END
  END OUT_IC_data[19]
  PIN OUT_IC_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2810.080 4.000 2810.640 ;
    END
  END OUT_IC_data[1]
  PIN OUT_IC_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2205.280 4.000 2205.840 ;
    END
  END OUT_IC_data[20]
  PIN OUT_IC_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2182.880 4.000 2183.440 ;
    END
  END OUT_IC_data[21]
  PIN OUT_IC_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2160.480 4.000 2161.040 ;
    END
  END OUT_IC_data[22]
  PIN OUT_IC_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2138.080 4.000 2138.640 ;
    END
  END OUT_IC_data[23]
  PIN OUT_IC_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2115.680 4.000 2116.240 ;
    END
  END OUT_IC_data[24]
  PIN OUT_IC_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2093.280 4.000 2093.840 ;
    END
  END OUT_IC_data[25]
  PIN OUT_IC_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2070.880 4.000 2071.440 ;
    END
  END OUT_IC_data[26]
  PIN OUT_IC_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2048.480 4.000 2049.040 ;
    END
  END OUT_IC_data[27]
  PIN OUT_IC_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2026.080 4.000 2026.640 ;
    END
  END OUT_IC_data[28]
  PIN OUT_IC_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2003.680 4.000 2004.240 ;
    END
  END OUT_IC_data[29]
  PIN OUT_IC_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2765.280 4.000 2765.840 ;
    END
  END OUT_IC_data[2]
  PIN OUT_IC_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1981.280 4.000 1981.840 ;
    END
  END OUT_IC_data[30]
  PIN OUT_IC_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1958.880 4.000 1959.440 ;
    END
  END OUT_IC_data[31]
  PIN OUT_IC_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2720.480 4.000 2721.040 ;
    END
  END OUT_IC_data[3]
  PIN OUT_IC_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2675.680 4.000 2676.240 ;
    END
  END OUT_IC_data[4]
  PIN OUT_IC_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2630.880 4.000 2631.440 ;
    END
  END OUT_IC_data[5]
  PIN OUT_IC_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2586.080 4.000 2586.640 ;
    END
  END OUT_IC_data[6]
  PIN OUT_IC_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2541.280 4.000 2541.840 ;
    END
  END OUT_IC_data[7]
  PIN OUT_IC_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2496.480 4.000 2497.040 ;
    END
  END OUT_IC_data[8]
  PIN OUT_IC_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2451.680 4.000 2452.240 ;
    END
  END OUT_IC_data[9]
  PIN OUT_IC_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.953000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2922.080 4.000 2922.640 ;
    END
  END OUT_IC_we
  PIN OUT_IC_wm
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2899.680 4.000 2900.240 ;
    END
  END OUT_IC_wm
  PIN OUT_dbgMemC[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2261.280 0.000 2261.840 4.000 ;
    END
  END OUT_dbgMemC[0]
  PIN OUT_dbgMemC[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2485.280 0.000 2485.840 4.000 ;
    END
  END OUT_dbgMemC[10]
  PIN OUT_dbgMemC[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2507.680 0.000 2508.240 4.000 ;
    END
  END OUT_dbgMemC[11]
  PIN OUT_dbgMemC[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.855000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2530.080 0.000 2530.640 4.000 ;
    END
  END OUT_dbgMemC[12]
  PIN OUT_dbgMemC[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.555500 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2552.480 0.000 2553.040 4.000 ;
    END
  END OUT_dbgMemC[13]
  PIN OUT_dbgMemC[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2574.880 0.000 2575.440 4.000 ;
    END
  END OUT_dbgMemC[14]
  PIN OUT_dbgMemC[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2597.280 0.000 2597.840 4.000 ;
    END
  END OUT_dbgMemC[15]
  PIN OUT_dbgMemC[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2283.680 0.000 2284.240 4.000 ;
    END
  END OUT_dbgMemC[1]
  PIN OUT_dbgMemC[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2306.080 0.000 2306.640 4.000 ;
    END
  END OUT_dbgMemC[2]
  PIN OUT_dbgMemC[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2328.480 0.000 2329.040 4.000 ;
    END
  END OUT_dbgMemC[3]
  PIN OUT_dbgMemC[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.261000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2350.880 0.000 2351.440 4.000 ;
    END
  END OUT_dbgMemC[4]
  PIN OUT_dbgMemC[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.261000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2373.280 0.000 2373.840 4.000 ;
    END
  END OUT_dbgMemC[5]
  PIN OUT_dbgMemC[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2395.680 0.000 2396.240 4.000 ;
    END
  END OUT_dbgMemC[6]
  PIN OUT_dbgMemC[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2418.080 0.000 2418.640 4.000 ;
    END
  END OUT_dbgMemC[7]
  PIN OUT_dbgMemC[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.804000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2440.480 0.000 2441.040 4.000 ;
    END
  END OUT_dbgMemC[8]
  PIN OUT_dbgMemC[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.002000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2462.880 0.000 2463.440 4.000 ;
    END
  END OUT_dbgMemC[9]
  PIN OUT_dbg[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2250.080 0.000 2250.640 4.000 ;
    END
  END OUT_dbg[0]
  PIN OUT_dbg[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2474.080 0.000 2474.640 4.000 ;
    END
  END OUT_dbg[10]
  PIN OUT_dbg[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2496.480 0.000 2497.040 4.000 ;
    END
  END OUT_dbg[11]
  PIN OUT_dbg[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2518.880 0.000 2519.440 4.000 ;
    END
  END OUT_dbg[12]
  PIN OUT_dbg[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2541.280 0.000 2541.840 4.000 ;
    END
  END OUT_dbg[13]
  PIN OUT_dbg[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2563.680 0.000 2564.240 4.000 ;
    END
  END OUT_dbg[14]
  PIN OUT_dbg[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2586.080 0.000 2586.640 4.000 ;
    END
  END OUT_dbg[15]
  PIN OUT_dbg[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2608.480 0.000 2609.040 4.000 ;
    END
  END OUT_dbg[16]
  PIN OUT_dbg[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2619.680 0.000 2620.240 4.000 ;
    END
  END OUT_dbg[17]
  PIN OUT_dbg[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2630.880 0.000 2631.440 4.000 ;
    END
  END OUT_dbg[18]
  PIN OUT_dbg[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2642.080 0.000 2642.640 4.000 ;
    END
  END OUT_dbg[19]
  PIN OUT_dbg[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2272.480 0.000 2273.040 4.000 ;
    END
  END OUT_dbg[1]
  PIN OUT_dbg[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2653.280 0.000 2653.840 4.000 ;
    END
  END OUT_dbg[20]
  PIN OUT_dbg[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2664.480 0.000 2665.040 4.000 ;
    END
  END OUT_dbg[21]
  PIN OUT_dbg[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2675.680 0.000 2676.240 4.000 ;
    END
  END OUT_dbg[22]
  PIN OUT_dbg[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2686.880 0.000 2687.440 4.000 ;
    END
  END OUT_dbg[23]
  PIN OUT_dbg[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2698.080 0.000 2698.640 4.000 ;
    END
  END OUT_dbg[24]
  PIN OUT_dbg[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2709.280 0.000 2709.840 4.000 ;
    END
  END OUT_dbg[25]
  PIN OUT_dbg[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2720.480 0.000 2721.040 4.000 ;
    END
  END OUT_dbg[26]
  PIN OUT_dbg[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2731.680 0.000 2732.240 4.000 ;
    END
  END OUT_dbg[27]
  PIN OUT_dbg[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2742.880 0.000 2743.440 4.000 ;
    END
  END OUT_dbg[28]
  PIN OUT_dbg[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2754.080 0.000 2754.640 4.000 ;
    END
  END OUT_dbg[29]
  PIN OUT_dbg[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2294.880 0.000 2295.440 4.000 ;
    END
  END OUT_dbg[2]
  PIN OUT_dbg[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2765.280 0.000 2765.840 4.000 ;
    END
  END OUT_dbg[30]
  PIN OUT_dbg[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2776.480 0.000 2777.040 4.000 ;
    END
  END OUT_dbg[31]
  PIN OUT_dbg[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2787.680 0.000 2788.240 4.000 ;
    END
  END OUT_dbg[32]
  PIN OUT_dbg[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2798.880 0.000 2799.440 4.000 ;
    END
  END OUT_dbg[33]
  PIN OUT_dbg[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2810.080 0.000 2810.640 4.000 ;
    END
  END OUT_dbg[34]
  PIN OUT_dbg[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2821.280 0.000 2821.840 4.000 ;
    END
  END OUT_dbg[35]
  PIN OUT_dbg[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2832.480 0.000 2833.040 4.000 ;
    END
  END OUT_dbg[36]
  PIN OUT_dbg[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2843.680 0.000 2844.240 4.000 ;
    END
  END OUT_dbg[37]
  PIN OUT_dbg[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2854.880 0.000 2855.440 4.000 ;
    END
  END OUT_dbg[38]
  PIN OUT_dbg[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2866.080 0.000 2866.640 4.000 ;
    END
  END OUT_dbg[39]
  PIN OUT_dbg[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.826000 ;
    ANTENNADIFFAREA 0.948400 ;
    PORT
      LAYER Metal2 ;
        RECT 2317.280 0.000 2317.840 4.000 ;
    END
  END OUT_dbg[3]
  PIN OUT_dbg[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.255500 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2339.680 0.000 2340.240 4.000 ;
    END
  END OUT_dbg[4]
  PIN OUT_dbg[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 1.672850 ;
    PORT
      LAYER Metal2 ;
        RECT 2362.080 0.000 2362.640 4.000 ;
    END
  END OUT_dbg[5]
  PIN OUT_dbg[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2384.480 0.000 2385.040 4.000 ;
    END
  END OUT_dbg[6]
  PIN OUT_dbg[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2406.880 0.000 2407.440 4.000 ;
    END
  END OUT_dbg[7]
  PIN OUT_dbg[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2429.280 0.000 2429.840 4.000 ;
    END
  END OUT_dbg[8]
  PIN OUT_dbg[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2451.680 0.000 2452.240 4.000 ;
    END
  END OUT_dbg[9]
  PIN OUT_powerOff
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2227.680 0.000 2228.240 4.000 ;
    END
  END OUT_powerOff
  PIN OUT_reboot
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2238.880 0.000 2239.440 4.000 ;
    END
  END OUT_reboot
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2194.080 0.000 2194.640 4.000 ;
    END
  END clk
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.914500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2216.480 0.000 2217.040 4.000 ;
    END
  END en
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.345500 ;
    ANTENNADIFFAREA 1.231200 ;
    PORT
      LAYER Metal2 ;
        RECT 2205.280 0.000 2205.840 4.000 ;
    END
  END rst
  PIN s_axi_araddr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 334.880 0.000 335.440 4.000 ;
    END
  END s_axi_araddr[0]
  PIN s_axi_araddr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1208.480 0.000 1209.040 4.000 ;
    END
  END s_axi_araddr[10]
  PIN s_axi_araddr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1253.280 0.000 1253.840 4.000 ;
    END
  END s_axi_araddr[11]
  PIN s_axi_araddr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1298.080 0.000 1298.640 4.000 ;
    END
  END s_axi_araddr[12]
  PIN s_axi_araddr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1342.880 0.000 1343.440 4.000 ;
    END
  END s_axi_araddr[13]
  PIN s_axi_araddr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1387.680 0.000 1388.240 4.000 ;
    END
  END s_axi_araddr[14]
  PIN s_axi_araddr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1432.480 0.000 1433.040 4.000 ;
    END
  END s_axi_araddr[15]
  PIN s_axi_araddr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1477.280 0.000 1477.840 4.000 ;
    END
  END s_axi_araddr[16]
  PIN s_axi_araddr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1522.080 0.000 1522.640 4.000 ;
    END
  END s_axi_araddr[17]
  PIN s_axi_araddr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1566.880 0.000 1567.440 4.000 ;
    END
  END s_axi_araddr[18]
  PIN s_axi_araddr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1611.680 0.000 1612.240 4.000 ;
    END
  END s_axi_araddr[19]
  PIN s_axi_araddr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 480.480 0.000 481.040 4.000 ;
    END
  END s_axi_araddr[1]
  PIN s_axi_araddr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1656.480 0.000 1657.040 4.000 ;
    END
  END s_axi_araddr[20]
  PIN s_axi_araddr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1701.280 0.000 1701.840 4.000 ;
    END
  END s_axi_araddr[21]
  PIN s_axi_araddr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1746.080 0.000 1746.640 4.000 ;
    END
  END s_axi_araddr[22]
  PIN s_axi_araddr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1790.880 0.000 1791.440 4.000 ;
    END
  END s_axi_araddr[23]
  PIN s_axi_araddr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1835.680 0.000 1836.240 4.000 ;
    END
  END s_axi_araddr[24]
  PIN s_axi_araddr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1880.480 0.000 1881.040 4.000 ;
    END
  END s_axi_araddr[25]
  PIN s_axi_araddr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1925.280 0.000 1925.840 4.000 ;
    END
  END s_axi_araddr[26]
  PIN s_axi_araddr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1970.080 0.000 1970.640 4.000 ;
    END
  END s_axi_araddr[27]
  PIN s_axi_araddr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 2014.880 0.000 2015.440 4.000 ;
    END
  END s_axi_araddr[28]
  PIN s_axi_araddr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 2059.680 0.000 2060.240 4.000 ;
    END
  END s_axi_araddr[29]
  PIN s_axi_araddr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 626.080 0.000 626.640 4.000 ;
    END
  END s_axi_araddr[2]
  PIN s_axi_araddr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 2104.480 0.000 2105.040 4.000 ;
    END
  END s_axi_araddr[30]
  PIN s_axi_araddr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 2149.280 0.000 2149.840 4.000 ;
    END
  END s_axi_araddr[31]
  PIN s_axi_araddr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 749.280 0.000 749.840 4.000 ;
    END
  END s_axi_araddr[3]
  PIN s_axi_araddr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 850.080 0.000 850.640 4.000 ;
    END
  END s_axi_araddr[4]
  PIN s_axi_araddr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 917.280 0.000 917.840 4.000 ;
    END
  END s_axi_araddr[5]
  PIN s_axi_araddr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 984.480 0.000 985.040 4.000 ;
    END
  END s_axi_araddr[6]
  PIN s_axi_araddr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1051.680 0.000 1052.240 4.000 ;
    END
  END s_axi_araddr[7]
  PIN s_axi_araddr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1118.880 0.000 1119.440 4.000 ;
    END
  END s_axi_araddr[8]
  PIN s_axi_araddr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1163.680 0.000 1164.240 4.000 ;
    END
  END s_axi_araddr[9]
  PIN s_axi_arburst[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 346.080 0.000 346.640 4.000 ;
    END
  END s_axi_arburst[0]
  PIN s_axi_arburst[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.997000 ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 491.680 0.000 492.240 4.000 ;
    END
  END s_axi_arburst[1]
  PIN s_axi_arcache[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 357.280 0.000 357.840 4.000 ;
    END
  END s_axi_arcache[0]
  PIN s_axi_arcache[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 502.880 0.000 503.440 4.000 ;
    END
  END s_axi_arcache[1]
  PIN s_axi_arcache[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 637.280 0.000 637.840 4.000 ;
    END
  END s_axi_arcache[2]
  PIN s_axi_arcache[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 760.480 0.000 761.040 4.000 ;
    END
  END s_axi_arcache[3]
  PIN s_axi_arid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 133.280 0.000 133.840 4.000 ;
    END
  END s_axi_arid
  PIN s_axi_arlen[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 368.480 0.000 369.040 4.000 ;
    END
  END s_axi_arlen[0]
  PIN s_axi_arlen[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 514.080 0.000 514.640 4.000 ;
    END
  END s_axi_arlen[1]
  PIN s_axi_arlen[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 648.480 0.000 649.040 4.000 ;
    END
  END s_axi_arlen[2]
  PIN s_axi_arlen[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 771.680 0.000 772.240 4.000 ;
    END
  END s_axi_arlen[3]
  PIN s_axi_arlen[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 861.280 0.000 861.840 4.000 ;
    END
  END s_axi_arlen[4]
  PIN s_axi_arlen[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 928.480 0.000 929.040 4.000 ;
    END
  END s_axi_arlen[5]
  PIN s_axi_arlen[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 995.680 0.000 996.240 4.000 ;
    END
  END s_axi_arlen[6]
  PIN s_axi_arlen[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1062.880 0.000 1063.440 4.000 ;
    END
  END s_axi_arlen[7]
  PIN s_axi_arlock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 0.000 145.040 4.000 ;
    END
  END s_axi_arlock
  PIN s_axi_arready
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.994500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 0.000 156.240 4.000 ;
    END
  END s_axi_arready
  PIN s_axi_arsize[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 379.680 0.000 380.240 4.000 ;
    END
  END s_axi_arsize[0]
  PIN s_axi_arsize[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 525.280 0.000 525.840 4.000 ;
    END
  END s_axi_arsize[1]
  PIN s_axi_arsize[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 659.680 0.000 660.240 4.000 ;
    END
  END s_axi_arsize[2]
  PIN s_axi_arvalid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 166.880 0.000 167.440 4.000 ;
    END
  END s_axi_arvalid
  PIN s_axi_awaddr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 390.880 0.000 391.440 4.000 ;
    END
  END s_axi_awaddr[0]
  PIN s_axi_awaddr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1219.680 0.000 1220.240 4.000 ;
    END
  END s_axi_awaddr[10]
  PIN s_axi_awaddr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1264.480 0.000 1265.040 4.000 ;
    END
  END s_axi_awaddr[11]
  PIN s_axi_awaddr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1309.280 0.000 1309.840 4.000 ;
    END
  END s_axi_awaddr[12]
  PIN s_axi_awaddr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1354.080 0.000 1354.640 4.000 ;
    END
  END s_axi_awaddr[13]
  PIN s_axi_awaddr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1398.880 0.000 1399.440 4.000 ;
    END
  END s_axi_awaddr[14]
  PIN s_axi_awaddr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1443.680 0.000 1444.240 4.000 ;
    END
  END s_axi_awaddr[15]
  PIN s_axi_awaddr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1488.480 0.000 1489.040 4.000 ;
    END
  END s_axi_awaddr[16]
  PIN s_axi_awaddr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1533.280 0.000 1533.840 4.000 ;
    END
  END s_axi_awaddr[17]
  PIN s_axi_awaddr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1578.080 0.000 1578.640 4.000 ;
    END
  END s_axi_awaddr[18]
  PIN s_axi_awaddr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1622.880 0.000 1623.440 4.000 ;
    END
  END s_axi_awaddr[19]
  PIN s_axi_awaddr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 536.480 0.000 537.040 4.000 ;
    END
  END s_axi_awaddr[1]
  PIN s_axi_awaddr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1667.680 0.000 1668.240 4.000 ;
    END
  END s_axi_awaddr[20]
  PIN s_axi_awaddr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1712.480 0.000 1713.040 4.000 ;
    END
  END s_axi_awaddr[21]
  PIN s_axi_awaddr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1757.280 0.000 1757.840 4.000 ;
    END
  END s_axi_awaddr[22]
  PIN s_axi_awaddr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1802.080 0.000 1802.640 4.000 ;
    END
  END s_axi_awaddr[23]
  PIN s_axi_awaddr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1846.880 0.000 1847.440 4.000 ;
    END
  END s_axi_awaddr[24]
  PIN s_axi_awaddr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1891.680 0.000 1892.240 4.000 ;
    END
  END s_axi_awaddr[25]
  PIN s_axi_awaddr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1936.480 0.000 1937.040 4.000 ;
    END
  END s_axi_awaddr[26]
  PIN s_axi_awaddr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1981.280 0.000 1981.840 4.000 ;
    END
  END s_axi_awaddr[27]
  PIN s_axi_awaddr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 2026.080 0.000 2026.640 4.000 ;
    END
  END s_axi_awaddr[28]
  PIN s_axi_awaddr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 2070.880 0.000 2071.440 4.000 ;
    END
  END s_axi_awaddr[29]
  PIN s_axi_awaddr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 670.880 0.000 671.440 4.000 ;
    END
  END s_axi_awaddr[2]
  PIN s_axi_awaddr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 2115.680 0.000 2116.240 4.000 ;
    END
  END s_axi_awaddr[30]
  PIN s_axi_awaddr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 2160.480 0.000 2161.040 4.000 ;
    END
  END s_axi_awaddr[31]
  PIN s_axi_awaddr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 782.880 0.000 783.440 4.000 ;
    END
  END s_axi_awaddr[3]
  PIN s_axi_awaddr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 872.480 0.000 873.040 4.000 ;
    END
  END s_axi_awaddr[4]
  PIN s_axi_awaddr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 939.680 0.000 940.240 4.000 ;
    END
  END s_axi_awaddr[5]
  PIN s_axi_awaddr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1006.880 0.000 1007.440 4.000 ;
    END
  END s_axi_awaddr[6]
  PIN s_axi_awaddr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1074.080 0.000 1074.640 4.000 ;
    END
  END s_axi_awaddr[7]
  PIN s_axi_awaddr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1130.080 0.000 1130.640 4.000 ;
    END
  END s_axi_awaddr[8]
  PIN s_axi_awaddr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 1174.880 0.000 1175.440 4.000 ;
    END
  END s_axi_awaddr[9]
  PIN s_axi_awburst[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 402.080 0.000 402.640 4.000 ;
    END
  END s_axi_awburst[0]
  PIN s_axi_awburst[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.997000 ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 547.680 0.000 548.240 4.000 ;
    END
  END s_axi_awburst[1]
  PIN s_axi_awcache[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 413.280 0.000 413.840 4.000 ;
    END
  END s_axi_awcache[0]
  PIN s_axi_awcache[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 558.880 0.000 559.440 4.000 ;
    END
  END s_axi_awcache[1]
  PIN s_axi_awcache[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 682.080 0.000 682.640 4.000 ;
    END
  END s_axi_awcache[2]
  PIN s_axi_awcache[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 794.080 0.000 794.640 4.000 ;
    END
  END s_axi_awcache[3]
  PIN s_axi_awid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 0.000 178.640 4.000 ;
    END
  END s_axi_awid
  PIN s_axi_awlen[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 424.480 0.000 425.040 4.000 ;
    END
  END s_axi_awlen[0]
  PIN s_axi_awlen[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 570.080 0.000 570.640 4.000 ;
    END
  END s_axi_awlen[1]
  PIN s_axi_awlen[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 693.280 0.000 693.840 4.000 ;
    END
  END s_axi_awlen[2]
  PIN s_axi_awlen[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 805.280 0.000 805.840 4.000 ;
    END
  END s_axi_awlen[3]
  PIN s_axi_awlen[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 883.680 0.000 884.240 4.000 ;
    END
  END s_axi_awlen[4]
  PIN s_axi_awlen[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 950.880 0.000 951.440 4.000 ;
    END
  END s_axi_awlen[5]
  PIN s_axi_awlen[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1018.080 0.000 1018.640 4.000 ;
    END
  END s_axi_awlen[6]
  PIN s_axi_awlen[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1085.280 0.000 1085.840 4.000 ;
    END
  END s_axi_awlen[7]
  PIN s_axi_awlock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 189.280 0.000 189.840 4.000 ;
    END
  END s_axi_awlock
  PIN s_axi_awready
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.994500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 200.480 0.000 201.040 4.000 ;
    END
  END s_axi_awready
  PIN s_axi_awsize[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 435.680 0.000 436.240 4.000 ;
    END
  END s_axi_awsize[0]
  PIN s_axi_awsize[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal2 ;
        RECT 581.280 0.000 581.840 4.000 ;
    END
  END s_axi_awsize[1]
  PIN s_axi_awsize[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 704.480 0.000 705.040 4.000 ;
    END
  END s_axi_awsize[2]
  PIN s_axi_awvalid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 0.000 212.240 4.000 ;
    END
  END s_axi_awvalid
  PIN s_axi_bid
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.092500 ;
    ANTENNADIFFAREA 1.641600 ;
    PORT
      LAYER Metal2 ;
        RECT 222.880 0.000 223.440 4.000 ;
    END
  END s_axi_bid
  PIN s_axi_bready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 234.080 0.000 234.640 4.000 ;
    END
  END s_axi_bready
  PIN s_axi_bvalid
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.576000 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 0.000 245.840 4.000 ;
    END
  END s_axi_bvalid
  PIN s_axi_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 446.880 0.000 447.440 4.000 ;
    END
  END s_axi_rdata[0]
  PIN s_axi_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 1230.880 0.000 1231.440 4.000 ;
    END
  END s_axi_rdata[10]
  PIN s_axi_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 1275.680 0.000 1276.240 4.000 ;
    END
  END s_axi_rdata[11]
  PIN s_axi_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 1320.480 0.000 1321.040 4.000 ;
    END
  END s_axi_rdata[12]
  PIN s_axi_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 1365.280 0.000 1365.840 4.000 ;
    END
  END s_axi_rdata[13]
  PIN s_axi_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 1410.080 0.000 1410.640 4.000 ;
    END
  END s_axi_rdata[14]
  PIN s_axi_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 1454.880 0.000 1455.440 4.000 ;
    END
  END s_axi_rdata[15]
  PIN s_axi_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 1499.680 0.000 1500.240 4.000 ;
    END
  END s_axi_rdata[16]
  PIN s_axi_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 1544.480 0.000 1545.040 4.000 ;
    END
  END s_axi_rdata[17]
  PIN s_axi_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 1589.280 0.000 1589.840 4.000 ;
    END
  END s_axi_rdata[18]
  PIN s_axi_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 1634.080 0.000 1634.640 4.000 ;
    END
  END s_axi_rdata[19]
  PIN s_axi_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 592.480 0.000 593.040 4.000 ;
    END
  END s_axi_rdata[1]
  PIN s_axi_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 1678.880 0.000 1679.440 4.000 ;
    END
  END s_axi_rdata[20]
  PIN s_axi_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 1723.680 0.000 1724.240 4.000 ;
    END
  END s_axi_rdata[21]
  PIN s_axi_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 1768.480 0.000 1769.040 4.000 ;
    END
  END s_axi_rdata[22]
  PIN s_axi_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 1813.280 0.000 1813.840 4.000 ;
    END
  END s_axi_rdata[23]
  PIN s_axi_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 1858.080 0.000 1858.640 4.000 ;
    END
  END s_axi_rdata[24]
  PIN s_axi_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 1902.880 0.000 1903.440 4.000 ;
    END
  END s_axi_rdata[25]
  PIN s_axi_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 1947.680 0.000 1948.240 4.000 ;
    END
  END s_axi_rdata[26]
  PIN s_axi_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 1992.480 0.000 1993.040 4.000 ;
    END
  END s_axi_rdata[27]
  PIN s_axi_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 2037.280 0.000 2037.840 4.000 ;
    END
  END s_axi_rdata[28]
  PIN s_axi_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 2082.080 0.000 2082.640 4.000 ;
    END
  END s_axi_rdata[29]
  PIN s_axi_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 715.680 0.000 716.240 4.000 ;
    END
  END s_axi_rdata[2]
  PIN s_axi_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 2126.880 0.000 2127.440 4.000 ;
    END
  END s_axi_rdata[30]
  PIN s_axi_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 2171.680 0.000 2172.240 4.000 ;
    END
  END s_axi_rdata[31]
  PIN s_axi_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 816.480 0.000 817.040 4.000 ;
    END
  END s_axi_rdata[3]
  PIN s_axi_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 894.880 0.000 895.440 4.000 ;
    END
  END s_axi_rdata[4]
  PIN s_axi_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 962.080 0.000 962.640 4.000 ;
    END
  END s_axi_rdata[5]
  PIN s_axi_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 1029.280 0.000 1029.840 4.000 ;
    END
  END s_axi_rdata[6]
  PIN s_axi_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 1096.480 0.000 1097.040 4.000 ;
    END
  END s_axi_rdata[7]
  PIN s_axi_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 1141.280 0.000 1141.840 4.000 ;
    END
  END s_axi_rdata[8]
  PIN s_axi_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.146500 ;
    ANTENNADIFFAREA 2.052000 ;
    PORT
      LAYER Metal2 ;
        RECT 1186.080 0.000 1186.640 4.000 ;
    END
  END s_axi_rdata[9]
  PIN s_axi_rid
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.997500 ;
    ANTENNADIFFAREA 0.820800 ;
    PORT
      LAYER Metal2 ;
        RECT 256.480 0.000 257.040 4.000 ;
    END
  END s_axi_rid
  PIN s_axi_rlast
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 267.680 0.000 268.240 4.000 ;
    END
  END s_axi_rlast
  PIN s_axi_rready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.984500 ;
    ANTENNADIFFAREA 1.306400 ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 0.000 279.440 4.000 ;
    END
  END s_axi_rready
  PIN s_axi_rvalid
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.041500 ;
    ANTENNADIFFAREA 1.641600 ;
    PORT
      LAYER Metal2 ;
        RECT 290.080 0.000 290.640 4.000 ;
    END
  END s_axi_rvalid
  PIN s_axi_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 458.080 0.000 458.640 4.000 ;
    END
  END s_axi_wdata[0]
  PIN s_axi_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1242.080 0.000 1242.640 4.000 ;
    END
  END s_axi_wdata[10]
  PIN s_axi_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1286.880 0.000 1287.440 4.000 ;
    END
  END s_axi_wdata[11]
  PIN s_axi_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1331.680 0.000 1332.240 4.000 ;
    END
  END s_axi_wdata[12]
  PIN s_axi_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1376.480 0.000 1377.040 4.000 ;
    END
  END s_axi_wdata[13]
  PIN s_axi_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1421.280 0.000 1421.840 4.000 ;
    END
  END s_axi_wdata[14]
  PIN s_axi_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1466.080 0.000 1466.640 4.000 ;
    END
  END s_axi_wdata[15]
  PIN s_axi_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1510.880 0.000 1511.440 4.000 ;
    END
  END s_axi_wdata[16]
  PIN s_axi_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1555.680 0.000 1556.240 4.000 ;
    END
  END s_axi_wdata[17]
  PIN s_axi_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1600.480 0.000 1601.040 4.000 ;
    END
  END s_axi_wdata[18]
  PIN s_axi_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1645.280 0.000 1645.840 4.000 ;
    END
  END s_axi_wdata[19]
  PIN s_axi_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 603.680 0.000 604.240 4.000 ;
    END
  END s_axi_wdata[1]
  PIN s_axi_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1690.080 0.000 1690.640 4.000 ;
    END
  END s_axi_wdata[20]
  PIN s_axi_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1734.880 0.000 1735.440 4.000 ;
    END
  END s_axi_wdata[21]
  PIN s_axi_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1779.680 0.000 1780.240 4.000 ;
    END
  END s_axi_wdata[22]
  PIN s_axi_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1824.480 0.000 1825.040 4.000 ;
    END
  END s_axi_wdata[23]
  PIN s_axi_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1869.280 0.000 1869.840 4.000 ;
    END
  END s_axi_wdata[24]
  PIN s_axi_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1914.080 0.000 1914.640 4.000 ;
    END
  END s_axi_wdata[25]
  PIN s_axi_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1958.880 0.000 1959.440 4.000 ;
    END
  END s_axi_wdata[26]
  PIN s_axi_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2003.680 0.000 2004.240 4.000 ;
    END
  END s_axi_wdata[27]
  PIN s_axi_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2048.480 0.000 2049.040 4.000 ;
    END
  END s_axi_wdata[28]
  PIN s_axi_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2093.280 0.000 2093.840 4.000 ;
    END
  END s_axi_wdata[29]
  PIN s_axi_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 726.880 0.000 727.440 4.000 ;
    END
  END s_axi_wdata[2]
  PIN s_axi_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2138.080 0.000 2138.640 4.000 ;
    END
  END s_axi_wdata[30]
  PIN s_axi_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 2182.880 0.000 2183.440 4.000 ;
    END
  END s_axi_wdata[31]
  PIN s_axi_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 827.680 0.000 828.240 4.000 ;
    END
  END s_axi_wdata[3]
  PIN s_axi_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 906.080 0.000 906.640 4.000 ;
    END
  END s_axi_wdata[4]
  PIN s_axi_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 973.280 0.000 973.840 4.000 ;
    END
  END s_axi_wdata[5]
  PIN s_axi_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1040.480 0.000 1041.040 4.000 ;
    END
  END s_axi_wdata[6]
  PIN s_axi_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1107.680 0.000 1108.240 4.000 ;
    END
  END s_axi_wdata[7]
  PIN s_axi_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1152.480 0.000 1153.040 4.000 ;
    END
  END s_axi_wdata[8]
  PIN s_axi_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1197.280 0.000 1197.840 4.000 ;
    END
  END s_axi_wdata[9]
  PIN s_axi_wlast
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.057000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 301.280 0.000 301.840 4.000 ;
    END
  END s_axi_wlast
  PIN s_axi_wready
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.949000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 312.480 0.000 313.040 4.000 ;
    END
  END s_axi_wready
  PIN s_axi_wstrb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 469.280 0.000 469.840 4.000 ;
    END
  END s_axi_wstrb[0]
  PIN s_axi_wstrb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 614.880 0.000 615.440 4.000 ;
    END
  END s_axi_wstrb[1]
  PIN s_axi_wstrb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 738.080 0.000 738.640 4.000 ;
    END
  END s_axi_wstrb[2]
  PIN s_axi_wstrb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 838.880 0.000 839.440 4.000 ;
    END
  END s_axi_wstrb[3]
  PIN s_axi_wvalid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 323.680 0.000 324.240 4.000 ;
    END
  END s_axi_wvalid
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1251.040 15.380 1252.640 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1404.640 15.380 1406.240 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1558.240 15.380 1559.840 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1711.840 15.380 1713.440 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1865.440 15.380 1867.040 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2019.040 15.380 2020.640 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2172.640 15.380 2174.240 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2326.240 15.380 2327.840 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2479.840 15.380 2481.440 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2633.440 15.380 2635.040 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2787.040 15.380 2788.640 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2940.640 15.380 2942.240 2983.420 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1327.840 15.380 1329.440 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1481.440 15.380 1483.040 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1635.040 15.380 1636.640 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1788.640 15.380 1790.240 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1942.240 15.380 1943.840 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2095.840 15.380 2097.440 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2249.440 15.380 2251.040 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2403.040 15.380 2404.640 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2556.640 15.380 2558.240 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2710.240 15.380 2711.840 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2863.840 15.380 2865.440 2983.420 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 14.710 2993.200 2985.770 ;
      LAYER Metal2 ;
        RECT 0.140 2995.700 20.980 2999.830 ;
        RECT 22.140 2995.700 43.380 2999.830 ;
        RECT 44.540 2995.700 65.780 2999.830 ;
        RECT 66.940 2995.700 88.180 2999.830 ;
        RECT 89.340 2995.700 110.580 2999.830 ;
        RECT 111.740 2995.700 132.980 2999.830 ;
        RECT 134.140 2995.700 155.380 2999.830 ;
        RECT 156.540 2995.700 177.780 2999.830 ;
        RECT 178.940 2995.700 200.180 2999.830 ;
        RECT 201.340 2995.700 222.580 2999.830 ;
        RECT 223.740 2995.700 244.980 2999.830 ;
        RECT 246.140 2995.700 267.380 2999.830 ;
        RECT 268.540 2995.700 289.780 2999.830 ;
        RECT 290.940 2995.700 312.180 2999.830 ;
        RECT 313.340 2995.700 334.580 2999.830 ;
        RECT 335.740 2995.700 356.980 2999.830 ;
        RECT 358.140 2995.700 379.380 2999.830 ;
        RECT 380.540 2995.700 401.780 2999.830 ;
        RECT 402.940 2995.700 424.180 2999.830 ;
        RECT 425.340 2995.700 446.580 2999.830 ;
        RECT 447.740 2995.700 468.980 2999.830 ;
        RECT 470.140 2995.700 491.380 2999.830 ;
        RECT 492.540 2995.700 513.780 2999.830 ;
        RECT 514.940 2995.700 536.180 2999.830 ;
        RECT 537.340 2995.700 558.580 2999.830 ;
        RECT 559.740 2995.700 580.980 2999.830 ;
        RECT 582.140 2995.700 603.380 2999.830 ;
        RECT 604.540 2995.700 625.780 2999.830 ;
        RECT 626.940 2995.700 648.180 2999.830 ;
        RECT 649.340 2995.700 670.580 2999.830 ;
        RECT 671.740 2995.700 692.980 2999.830 ;
        RECT 694.140 2995.700 715.380 2999.830 ;
        RECT 716.540 2995.700 737.780 2999.830 ;
        RECT 738.940 2995.700 760.180 2999.830 ;
        RECT 761.340 2995.700 782.580 2999.830 ;
        RECT 783.740 2995.700 804.980 2999.830 ;
        RECT 806.140 2995.700 827.380 2999.830 ;
        RECT 828.540 2995.700 849.780 2999.830 ;
        RECT 850.940 2995.700 872.180 2999.830 ;
        RECT 873.340 2995.700 894.580 2999.830 ;
        RECT 895.740 2995.700 916.980 2999.830 ;
        RECT 918.140 2995.700 939.380 2999.830 ;
        RECT 940.540 2995.700 961.780 2999.830 ;
        RECT 962.940 2995.700 984.180 2999.830 ;
        RECT 985.340 2995.700 1006.580 2999.830 ;
        RECT 1007.740 2995.700 1028.980 2999.830 ;
        RECT 1030.140 2995.700 1051.380 2999.830 ;
        RECT 1052.540 2995.700 1073.780 2999.830 ;
        RECT 1074.940 2995.700 1096.180 2999.830 ;
        RECT 1097.340 2995.700 1118.580 2999.830 ;
        RECT 1119.740 2995.700 1140.980 2999.830 ;
        RECT 1142.140 2995.700 1163.380 2999.830 ;
        RECT 1164.540 2995.700 1185.780 2999.830 ;
        RECT 1186.940 2995.700 1208.180 2999.830 ;
        RECT 1209.340 2995.700 1230.580 2999.830 ;
        RECT 1231.740 2995.700 1252.980 2999.830 ;
        RECT 1254.140 2995.700 1275.380 2999.830 ;
        RECT 1276.540 2995.700 1297.780 2999.830 ;
        RECT 1298.940 2995.700 1320.180 2999.830 ;
        RECT 1321.340 2995.700 1342.580 2999.830 ;
        RECT 1343.740 2995.700 1364.980 2999.830 ;
        RECT 1366.140 2995.700 1387.380 2999.830 ;
        RECT 1388.540 2995.700 1409.780 2999.830 ;
        RECT 1410.940 2995.700 1432.180 2999.830 ;
        RECT 1433.340 2995.700 1454.580 2999.830 ;
        RECT 1455.740 2995.700 1476.980 2999.830 ;
        RECT 1478.140 2995.700 1499.380 2999.830 ;
        RECT 1500.540 2995.700 1521.780 2999.830 ;
        RECT 1522.940 2995.700 1544.180 2999.830 ;
        RECT 1545.340 2995.700 1566.580 2999.830 ;
        RECT 1567.740 2995.700 1588.980 2999.830 ;
        RECT 1590.140 2995.700 1611.380 2999.830 ;
        RECT 1612.540 2995.700 1633.780 2999.830 ;
        RECT 1634.940 2995.700 1656.180 2999.830 ;
        RECT 1657.340 2995.700 1678.580 2999.830 ;
        RECT 1679.740 2995.700 1700.980 2999.830 ;
        RECT 1702.140 2995.700 1723.380 2999.830 ;
        RECT 1724.540 2995.700 1745.780 2999.830 ;
        RECT 1746.940 2995.700 1768.180 2999.830 ;
        RECT 1769.340 2995.700 1790.580 2999.830 ;
        RECT 1791.740 2995.700 1812.980 2999.830 ;
        RECT 1814.140 2995.700 1835.380 2999.830 ;
        RECT 1836.540 2995.700 1857.780 2999.830 ;
        RECT 1858.940 2995.700 1880.180 2999.830 ;
        RECT 1881.340 2995.700 1902.580 2999.830 ;
        RECT 1903.740 2995.700 1924.980 2999.830 ;
        RECT 1926.140 2995.700 1947.380 2999.830 ;
        RECT 1948.540 2995.700 1969.780 2999.830 ;
        RECT 1970.940 2995.700 1992.180 2999.830 ;
        RECT 1993.340 2995.700 2014.580 2999.830 ;
        RECT 2015.740 2995.700 2036.980 2999.830 ;
        RECT 2038.140 2995.700 2059.380 2999.830 ;
        RECT 2060.540 2995.700 2081.780 2999.830 ;
        RECT 2082.940 2995.700 2104.180 2999.830 ;
        RECT 2105.340 2995.700 2126.580 2999.830 ;
        RECT 2127.740 2995.700 2148.980 2999.830 ;
        RECT 2150.140 2995.700 2171.380 2999.830 ;
        RECT 2172.540 2995.700 2193.780 2999.830 ;
        RECT 2194.940 2995.700 2216.180 2999.830 ;
        RECT 2217.340 2995.700 2238.580 2999.830 ;
        RECT 2239.740 2995.700 2260.980 2999.830 ;
        RECT 2262.140 2995.700 2283.380 2999.830 ;
        RECT 2284.540 2995.700 2305.780 2999.830 ;
        RECT 2306.940 2995.700 2328.180 2999.830 ;
        RECT 2329.340 2995.700 2350.580 2999.830 ;
        RECT 2351.740 2995.700 2372.980 2999.830 ;
        RECT 2374.140 2995.700 2395.380 2999.830 ;
        RECT 2396.540 2995.700 2417.780 2999.830 ;
        RECT 2418.940 2995.700 2440.180 2999.830 ;
        RECT 2441.340 2995.700 2462.580 2999.830 ;
        RECT 2463.740 2995.700 2484.980 2999.830 ;
        RECT 2486.140 2995.700 2507.380 2999.830 ;
        RECT 2508.540 2995.700 2529.780 2999.830 ;
        RECT 2530.940 2995.700 2552.180 2999.830 ;
        RECT 2553.340 2995.700 2574.580 2999.830 ;
        RECT 2575.740 2995.700 2596.980 2999.830 ;
        RECT 2598.140 2995.700 2619.380 2999.830 ;
        RECT 2620.540 2995.700 2641.780 2999.830 ;
        RECT 2642.940 2995.700 2664.180 2999.830 ;
        RECT 2665.340 2995.700 2686.580 2999.830 ;
        RECT 2687.740 2995.700 2708.980 2999.830 ;
        RECT 2710.140 2995.700 2731.380 2999.830 ;
        RECT 2732.540 2995.700 2753.780 2999.830 ;
        RECT 2754.940 2995.700 2776.180 2999.830 ;
        RECT 2777.340 2995.700 2798.580 2999.830 ;
        RECT 2799.740 2995.700 2820.980 2999.830 ;
        RECT 2822.140 2995.700 2843.380 2999.830 ;
        RECT 2844.540 2995.700 2865.780 2999.830 ;
        RECT 2866.940 2995.700 2888.180 2999.830 ;
        RECT 2889.340 2995.700 2910.580 2999.830 ;
        RECT 2911.740 2995.700 2932.980 2999.830 ;
        RECT 2934.140 2995.700 2955.380 2999.830 ;
        RECT 2956.540 2995.700 2977.780 2999.830 ;
        RECT 2978.940 2995.700 2993.620 2999.830 ;
        RECT 0.140 4.300 2993.620 2995.700 ;
        RECT 0.140 0.090 132.980 4.300 ;
        RECT 134.140 0.090 144.180 4.300 ;
        RECT 145.340 0.090 155.380 4.300 ;
        RECT 156.540 0.090 166.580 4.300 ;
        RECT 167.740 0.090 177.780 4.300 ;
        RECT 178.940 0.090 188.980 4.300 ;
        RECT 190.140 0.090 200.180 4.300 ;
        RECT 201.340 0.090 211.380 4.300 ;
        RECT 212.540 0.090 222.580 4.300 ;
        RECT 223.740 0.090 233.780 4.300 ;
        RECT 234.940 0.090 244.980 4.300 ;
        RECT 246.140 0.090 256.180 4.300 ;
        RECT 257.340 0.090 267.380 4.300 ;
        RECT 268.540 0.090 278.580 4.300 ;
        RECT 279.740 0.090 289.780 4.300 ;
        RECT 290.940 0.090 300.980 4.300 ;
        RECT 302.140 0.090 312.180 4.300 ;
        RECT 313.340 0.090 323.380 4.300 ;
        RECT 324.540 0.090 334.580 4.300 ;
        RECT 335.740 0.090 345.780 4.300 ;
        RECT 346.940 0.090 356.980 4.300 ;
        RECT 358.140 0.090 368.180 4.300 ;
        RECT 369.340 0.090 379.380 4.300 ;
        RECT 380.540 0.090 390.580 4.300 ;
        RECT 391.740 0.090 401.780 4.300 ;
        RECT 402.940 0.090 412.980 4.300 ;
        RECT 414.140 0.090 424.180 4.300 ;
        RECT 425.340 0.090 435.380 4.300 ;
        RECT 436.540 0.090 446.580 4.300 ;
        RECT 447.740 0.090 457.780 4.300 ;
        RECT 458.940 0.090 468.980 4.300 ;
        RECT 470.140 0.090 480.180 4.300 ;
        RECT 481.340 0.090 491.380 4.300 ;
        RECT 492.540 0.090 502.580 4.300 ;
        RECT 503.740 0.090 513.780 4.300 ;
        RECT 514.940 0.090 524.980 4.300 ;
        RECT 526.140 0.090 536.180 4.300 ;
        RECT 537.340 0.090 547.380 4.300 ;
        RECT 548.540 0.090 558.580 4.300 ;
        RECT 559.740 0.090 569.780 4.300 ;
        RECT 570.940 0.090 580.980 4.300 ;
        RECT 582.140 0.090 592.180 4.300 ;
        RECT 593.340 0.090 603.380 4.300 ;
        RECT 604.540 0.090 614.580 4.300 ;
        RECT 615.740 0.090 625.780 4.300 ;
        RECT 626.940 0.090 636.980 4.300 ;
        RECT 638.140 0.090 648.180 4.300 ;
        RECT 649.340 0.090 659.380 4.300 ;
        RECT 660.540 0.090 670.580 4.300 ;
        RECT 671.740 0.090 681.780 4.300 ;
        RECT 682.940 0.090 692.980 4.300 ;
        RECT 694.140 0.090 704.180 4.300 ;
        RECT 705.340 0.090 715.380 4.300 ;
        RECT 716.540 0.090 726.580 4.300 ;
        RECT 727.740 0.090 737.780 4.300 ;
        RECT 738.940 0.090 748.980 4.300 ;
        RECT 750.140 0.090 760.180 4.300 ;
        RECT 761.340 0.090 771.380 4.300 ;
        RECT 772.540 0.090 782.580 4.300 ;
        RECT 783.740 0.090 793.780 4.300 ;
        RECT 794.940 0.090 804.980 4.300 ;
        RECT 806.140 0.090 816.180 4.300 ;
        RECT 817.340 0.090 827.380 4.300 ;
        RECT 828.540 0.090 838.580 4.300 ;
        RECT 839.740 0.090 849.780 4.300 ;
        RECT 850.940 0.090 860.980 4.300 ;
        RECT 862.140 0.090 872.180 4.300 ;
        RECT 873.340 0.090 883.380 4.300 ;
        RECT 884.540 0.090 894.580 4.300 ;
        RECT 895.740 0.090 905.780 4.300 ;
        RECT 906.940 0.090 916.980 4.300 ;
        RECT 918.140 0.090 928.180 4.300 ;
        RECT 929.340 0.090 939.380 4.300 ;
        RECT 940.540 0.090 950.580 4.300 ;
        RECT 951.740 0.090 961.780 4.300 ;
        RECT 962.940 0.090 972.980 4.300 ;
        RECT 974.140 0.090 984.180 4.300 ;
        RECT 985.340 0.090 995.380 4.300 ;
        RECT 996.540 0.090 1006.580 4.300 ;
        RECT 1007.740 0.090 1017.780 4.300 ;
        RECT 1018.940 0.090 1028.980 4.300 ;
        RECT 1030.140 0.090 1040.180 4.300 ;
        RECT 1041.340 0.090 1051.380 4.300 ;
        RECT 1052.540 0.090 1062.580 4.300 ;
        RECT 1063.740 0.090 1073.780 4.300 ;
        RECT 1074.940 0.090 1084.980 4.300 ;
        RECT 1086.140 0.090 1096.180 4.300 ;
        RECT 1097.340 0.090 1107.380 4.300 ;
        RECT 1108.540 0.090 1118.580 4.300 ;
        RECT 1119.740 0.090 1129.780 4.300 ;
        RECT 1130.940 0.090 1140.980 4.300 ;
        RECT 1142.140 0.090 1152.180 4.300 ;
        RECT 1153.340 0.090 1163.380 4.300 ;
        RECT 1164.540 0.090 1174.580 4.300 ;
        RECT 1175.740 0.090 1185.780 4.300 ;
        RECT 1186.940 0.090 1196.980 4.300 ;
        RECT 1198.140 0.090 1208.180 4.300 ;
        RECT 1209.340 0.090 1219.380 4.300 ;
        RECT 1220.540 0.090 1230.580 4.300 ;
        RECT 1231.740 0.090 1241.780 4.300 ;
        RECT 1242.940 0.090 1252.980 4.300 ;
        RECT 1254.140 0.090 1264.180 4.300 ;
        RECT 1265.340 0.090 1275.380 4.300 ;
        RECT 1276.540 0.090 1286.580 4.300 ;
        RECT 1287.740 0.090 1297.780 4.300 ;
        RECT 1298.940 0.090 1308.980 4.300 ;
        RECT 1310.140 0.090 1320.180 4.300 ;
        RECT 1321.340 0.090 1331.380 4.300 ;
        RECT 1332.540 0.090 1342.580 4.300 ;
        RECT 1343.740 0.090 1353.780 4.300 ;
        RECT 1354.940 0.090 1364.980 4.300 ;
        RECT 1366.140 0.090 1376.180 4.300 ;
        RECT 1377.340 0.090 1387.380 4.300 ;
        RECT 1388.540 0.090 1398.580 4.300 ;
        RECT 1399.740 0.090 1409.780 4.300 ;
        RECT 1410.940 0.090 1420.980 4.300 ;
        RECT 1422.140 0.090 1432.180 4.300 ;
        RECT 1433.340 0.090 1443.380 4.300 ;
        RECT 1444.540 0.090 1454.580 4.300 ;
        RECT 1455.740 0.090 1465.780 4.300 ;
        RECT 1466.940 0.090 1476.980 4.300 ;
        RECT 1478.140 0.090 1488.180 4.300 ;
        RECT 1489.340 0.090 1499.380 4.300 ;
        RECT 1500.540 0.090 1510.580 4.300 ;
        RECT 1511.740 0.090 1521.780 4.300 ;
        RECT 1522.940 0.090 1532.980 4.300 ;
        RECT 1534.140 0.090 1544.180 4.300 ;
        RECT 1545.340 0.090 1555.380 4.300 ;
        RECT 1556.540 0.090 1566.580 4.300 ;
        RECT 1567.740 0.090 1577.780 4.300 ;
        RECT 1578.940 0.090 1588.980 4.300 ;
        RECT 1590.140 0.090 1600.180 4.300 ;
        RECT 1601.340 0.090 1611.380 4.300 ;
        RECT 1612.540 0.090 1622.580 4.300 ;
        RECT 1623.740 0.090 1633.780 4.300 ;
        RECT 1634.940 0.090 1644.980 4.300 ;
        RECT 1646.140 0.090 1656.180 4.300 ;
        RECT 1657.340 0.090 1667.380 4.300 ;
        RECT 1668.540 0.090 1678.580 4.300 ;
        RECT 1679.740 0.090 1689.780 4.300 ;
        RECT 1690.940 0.090 1700.980 4.300 ;
        RECT 1702.140 0.090 1712.180 4.300 ;
        RECT 1713.340 0.090 1723.380 4.300 ;
        RECT 1724.540 0.090 1734.580 4.300 ;
        RECT 1735.740 0.090 1745.780 4.300 ;
        RECT 1746.940 0.090 1756.980 4.300 ;
        RECT 1758.140 0.090 1768.180 4.300 ;
        RECT 1769.340 0.090 1779.380 4.300 ;
        RECT 1780.540 0.090 1790.580 4.300 ;
        RECT 1791.740 0.090 1801.780 4.300 ;
        RECT 1802.940 0.090 1812.980 4.300 ;
        RECT 1814.140 0.090 1824.180 4.300 ;
        RECT 1825.340 0.090 1835.380 4.300 ;
        RECT 1836.540 0.090 1846.580 4.300 ;
        RECT 1847.740 0.090 1857.780 4.300 ;
        RECT 1858.940 0.090 1868.980 4.300 ;
        RECT 1870.140 0.090 1880.180 4.300 ;
        RECT 1881.340 0.090 1891.380 4.300 ;
        RECT 1892.540 0.090 1902.580 4.300 ;
        RECT 1903.740 0.090 1913.780 4.300 ;
        RECT 1914.940 0.090 1924.980 4.300 ;
        RECT 1926.140 0.090 1936.180 4.300 ;
        RECT 1937.340 0.090 1947.380 4.300 ;
        RECT 1948.540 0.090 1958.580 4.300 ;
        RECT 1959.740 0.090 1969.780 4.300 ;
        RECT 1970.940 0.090 1980.980 4.300 ;
        RECT 1982.140 0.090 1992.180 4.300 ;
        RECT 1993.340 0.090 2003.380 4.300 ;
        RECT 2004.540 0.090 2014.580 4.300 ;
        RECT 2015.740 0.090 2025.780 4.300 ;
        RECT 2026.940 0.090 2036.980 4.300 ;
        RECT 2038.140 0.090 2048.180 4.300 ;
        RECT 2049.340 0.090 2059.380 4.300 ;
        RECT 2060.540 0.090 2070.580 4.300 ;
        RECT 2071.740 0.090 2081.780 4.300 ;
        RECT 2082.940 0.090 2092.980 4.300 ;
        RECT 2094.140 0.090 2104.180 4.300 ;
        RECT 2105.340 0.090 2115.380 4.300 ;
        RECT 2116.540 0.090 2126.580 4.300 ;
        RECT 2127.740 0.090 2137.780 4.300 ;
        RECT 2138.940 0.090 2148.980 4.300 ;
        RECT 2150.140 0.090 2160.180 4.300 ;
        RECT 2161.340 0.090 2171.380 4.300 ;
        RECT 2172.540 0.090 2182.580 4.300 ;
        RECT 2183.740 0.090 2193.780 4.300 ;
        RECT 2194.940 0.090 2204.980 4.300 ;
        RECT 2206.140 0.090 2216.180 4.300 ;
        RECT 2217.340 0.090 2227.380 4.300 ;
        RECT 2228.540 0.090 2238.580 4.300 ;
        RECT 2239.740 0.090 2249.780 4.300 ;
        RECT 2250.940 0.090 2260.980 4.300 ;
        RECT 2262.140 0.090 2272.180 4.300 ;
        RECT 2273.340 0.090 2283.380 4.300 ;
        RECT 2284.540 0.090 2294.580 4.300 ;
        RECT 2295.740 0.090 2305.780 4.300 ;
        RECT 2306.940 0.090 2316.980 4.300 ;
        RECT 2318.140 0.090 2328.180 4.300 ;
        RECT 2329.340 0.090 2339.380 4.300 ;
        RECT 2340.540 0.090 2350.580 4.300 ;
        RECT 2351.740 0.090 2361.780 4.300 ;
        RECT 2362.940 0.090 2372.980 4.300 ;
        RECT 2374.140 0.090 2384.180 4.300 ;
        RECT 2385.340 0.090 2395.380 4.300 ;
        RECT 2396.540 0.090 2406.580 4.300 ;
        RECT 2407.740 0.090 2417.780 4.300 ;
        RECT 2418.940 0.090 2428.980 4.300 ;
        RECT 2430.140 0.090 2440.180 4.300 ;
        RECT 2441.340 0.090 2451.380 4.300 ;
        RECT 2452.540 0.090 2462.580 4.300 ;
        RECT 2463.740 0.090 2473.780 4.300 ;
        RECT 2474.940 0.090 2484.980 4.300 ;
        RECT 2486.140 0.090 2496.180 4.300 ;
        RECT 2497.340 0.090 2507.380 4.300 ;
        RECT 2508.540 0.090 2518.580 4.300 ;
        RECT 2519.740 0.090 2529.780 4.300 ;
        RECT 2530.940 0.090 2540.980 4.300 ;
        RECT 2542.140 0.090 2552.180 4.300 ;
        RECT 2553.340 0.090 2563.380 4.300 ;
        RECT 2564.540 0.090 2574.580 4.300 ;
        RECT 2575.740 0.090 2585.780 4.300 ;
        RECT 2586.940 0.090 2596.980 4.300 ;
        RECT 2598.140 0.090 2608.180 4.300 ;
        RECT 2609.340 0.090 2619.380 4.300 ;
        RECT 2620.540 0.090 2630.580 4.300 ;
        RECT 2631.740 0.090 2641.780 4.300 ;
        RECT 2642.940 0.090 2652.980 4.300 ;
        RECT 2654.140 0.090 2664.180 4.300 ;
        RECT 2665.340 0.090 2675.380 4.300 ;
        RECT 2676.540 0.090 2686.580 4.300 ;
        RECT 2687.740 0.090 2697.780 4.300 ;
        RECT 2698.940 0.090 2708.980 4.300 ;
        RECT 2710.140 0.090 2720.180 4.300 ;
        RECT 2721.340 0.090 2731.380 4.300 ;
        RECT 2732.540 0.090 2742.580 4.300 ;
        RECT 2743.740 0.090 2753.780 4.300 ;
        RECT 2754.940 0.090 2764.980 4.300 ;
        RECT 2766.140 0.090 2776.180 4.300 ;
        RECT 2777.340 0.090 2787.380 4.300 ;
        RECT 2788.540 0.090 2798.580 4.300 ;
        RECT 2799.740 0.090 2809.780 4.300 ;
        RECT 2810.940 0.090 2820.980 4.300 ;
        RECT 2822.140 0.090 2832.180 4.300 ;
        RECT 2833.340 0.090 2843.380 4.300 ;
        RECT 2844.540 0.090 2854.580 4.300 ;
        RECT 2855.740 0.090 2865.780 4.300 ;
        RECT 2866.940 0.090 2993.620 4.300 ;
      LAYER Metal3 ;
        RECT 0.090 2945.340 2993.670 2999.780 ;
        RECT 4.300 2944.180 2993.670 2945.340 ;
        RECT 0.090 2922.940 2993.670 2944.180 ;
        RECT 4.300 2921.780 2993.670 2922.940 ;
        RECT 0.090 2900.540 2993.670 2921.780 ;
        RECT 4.300 2899.380 2993.670 2900.540 ;
        RECT 0.090 2878.140 2993.670 2899.380 ;
        RECT 4.300 2876.980 2993.670 2878.140 ;
        RECT 0.090 2855.740 2993.670 2876.980 ;
        RECT 4.300 2854.580 2993.670 2855.740 ;
        RECT 0.090 2833.340 2993.670 2854.580 ;
        RECT 4.300 2832.180 2993.670 2833.340 ;
        RECT 0.090 2810.940 2993.670 2832.180 ;
        RECT 4.300 2809.780 2993.670 2810.940 ;
        RECT 0.090 2788.540 2993.670 2809.780 ;
        RECT 4.300 2787.380 2993.670 2788.540 ;
        RECT 0.090 2766.140 2993.670 2787.380 ;
        RECT 4.300 2764.980 2993.670 2766.140 ;
        RECT 0.090 2743.740 2993.670 2764.980 ;
        RECT 4.300 2742.580 2993.670 2743.740 ;
        RECT 0.090 2721.340 2993.670 2742.580 ;
        RECT 4.300 2720.180 2993.670 2721.340 ;
        RECT 0.090 2698.940 2993.670 2720.180 ;
        RECT 4.300 2697.780 2993.670 2698.940 ;
        RECT 0.090 2676.540 2993.670 2697.780 ;
        RECT 4.300 2675.380 2993.670 2676.540 ;
        RECT 0.090 2654.140 2993.670 2675.380 ;
        RECT 4.300 2652.980 2993.670 2654.140 ;
        RECT 0.090 2631.740 2993.670 2652.980 ;
        RECT 4.300 2630.580 2993.670 2631.740 ;
        RECT 0.090 2609.340 2993.670 2630.580 ;
        RECT 4.300 2608.180 2993.670 2609.340 ;
        RECT 0.090 2586.940 2993.670 2608.180 ;
        RECT 4.300 2585.780 2993.670 2586.940 ;
        RECT 0.090 2564.540 2993.670 2585.780 ;
        RECT 4.300 2563.380 2993.670 2564.540 ;
        RECT 0.090 2542.140 2993.670 2563.380 ;
        RECT 4.300 2540.980 2993.670 2542.140 ;
        RECT 0.090 2519.740 2993.670 2540.980 ;
        RECT 4.300 2518.580 2993.670 2519.740 ;
        RECT 0.090 2497.340 2993.670 2518.580 ;
        RECT 4.300 2496.180 2993.670 2497.340 ;
        RECT 0.090 2474.940 2993.670 2496.180 ;
        RECT 4.300 2473.780 2993.670 2474.940 ;
        RECT 0.090 2452.540 2993.670 2473.780 ;
        RECT 4.300 2451.380 2993.670 2452.540 ;
        RECT 0.090 2430.140 2993.670 2451.380 ;
        RECT 4.300 2428.980 2993.670 2430.140 ;
        RECT 0.090 2407.740 2993.670 2428.980 ;
        RECT 4.300 2406.580 2993.670 2407.740 ;
        RECT 0.090 2385.340 2993.670 2406.580 ;
        RECT 4.300 2384.180 2993.670 2385.340 ;
        RECT 0.090 2362.940 2993.670 2384.180 ;
        RECT 4.300 2361.780 2993.670 2362.940 ;
        RECT 0.090 2340.540 2993.670 2361.780 ;
        RECT 4.300 2339.380 2993.670 2340.540 ;
        RECT 0.090 2318.140 2993.670 2339.380 ;
        RECT 4.300 2316.980 2993.670 2318.140 ;
        RECT 0.090 2295.740 2993.670 2316.980 ;
        RECT 4.300 2294.580 2993.670 2295.740 ;
        RECT 0.090 2273.340 2993.670 2294.580 ;
        RECT 4.300 2272.180 2993.670 2273.340 ;
        RECT 0.090 2250.940 2993.670 2272.180 ;
        RECT 4.300 2249.780 2993.670 2250.940 ;
        RECT 0.090 2228.540 2993.670 2249.780 ;
        RECT 4.300 2227.380 2993.670 2228.540 ;
        RECT 0.090 2206.140 2993.670 2227.380 ;
        RECT 4.300 2204.980 2993.670 2206.140 ;
        RECT 0.090 2183.740 2993.670 2204.980 ;
        RECT 4.300 2182.580 2993.670 2183.740 ;
        RECT 0.090 2161.340 2993.670 2182.580 ;
        RECT 4.300 2160.180 2993.670 2161.340 ;
        RECT 0.090 2138.940 2993.670 2160.180 ;
        RECT 4.300 2137.780 2993.670 2138.940 ;
        RECT 0.090 2116.540 2993.670 2137.780 ;
        RECT 4.300 2115.380 2993.670 2116.540 ;
        RECT 0.090 2094.140 2993.670 2115.380 ;
        RECT 4.300 2092.980 2993.670 2094.140 ;
        RECT 0.090 2071.740 2993.670 2092.980 ;
        RECT 4.300 2070.580 2993.670 2071.740 ;
        RECT 0.090 2049.340 2993.670 2070.580 ;
        RECT 4.300 2048.180 2993.670 2049.340 ;
        RECT 0.090 2026.940 2993.670 2048.180 ;
        RECT 4.300 2025.780 2993.670 2026.940 ;
        RECT 0.090 2004.540 2993.670 2025.780 ;
        RECT 4.300 2003.380 2993.670 2004.540 ;
        RECT 0.090 1982.140 2993.670 2003.380 ;
        RECT 4.300 1980.980 2993.670 1982.140 ;
        RECT 0.090 1959.740 2993.670 1980.980 ;
        RECT 4.300 1958.580 2993.670 1959.740 ;
        RECT 0.090 1937.340 2993.670 1958.580 ;
        RECT 4.300 1936.180 2993.670 1937.340 ;
        RECT 0.090 1914.940 2993.670 1936.180 ;
        RECT 4.300 1913.780 2993.670 1914.940 ;
        RECT 0.090 1892.540 2993.670 1913.780 ;
        RECT 4.300 1891.380 2993.670 1892.540 ;
        RECT 0.090 1870.140 2993.670 1891.380 ;
        RECT 4.300 1868.980 2993.670 1870.140 ;
        RECT 0.090 1847.740 2993.670 1868.980 ;
        RECT 4.300 1846.580 2993.670 1847.740 ;
        RECT 0.090 1825.340 2993.670 1846.580 ;
        RECT 4.300 1824.180 2993.670 1825.340 ;
        RECT 0.090 1802.940 2993.670 1824.180 ;
        RECT 4.300 1801.780 2993.670 1802.940 ;
        RECT 0.090 1780.540 2993.670 1801.780 ;
        RECT 4.300 1779.380 2993.670 1780.540 ;
        RECT 0.090 1758.140 2993.670 1779.380 ;
        RECT 4.300 1756.980 2993.670 1758.140 ;
        RECT 0.090 1735.740 2993.670 1756.980 ;
        RECT 4.300 1734.580 2993.670 1735.740 ;
        RECT 0.090 1713.340 2993.670 1734.580 ;
        RECT 4.300 1712.180 2993.670 1713.340 ;
        RECT 0.090 1690.940 2993.670 1712.180 ;
        RECT 4.300 1689.780 2993.670 1690.940 ;
        RECT 0.090 1668.540 2993.670 1689.780 ;
        RECT 4.300 1667.380 2993.670 1668.540 ;
        RECT 0.090 1646.140 2993.670 1667.380 ;
        RECT 4.300 1644.980 2993.670 1646.140 ;
        RECT 0.090 1623.740 2993.670 1644.980 ;
        RECT 4.300 1622.580 2993.670 1623.740 ;
        RECT 0.090 1601.340 2993.670 1622.580 ;
        RECT 4.300 1600.180 2993.670 1601.340 ;
        RECT 0.090 1578.940 2993.670 1600.180 ;
        RECT 4.300 1577.780 2993.670 1578.940 ;
        RECT 0.090 1556.540 2993.670 1577.780 ;
        RECT 4.300 1555.380 2993.670 1556.540 ;
        RECT 0.090 1534.140 2993.670 1555.380 ;
        RECT 4.300 1532.980 2993.670 1534.140 ;
        RECT 0.090 1511.740 2993.670 1532.980 ;
        RECT 4.300 1510.580 2993.670 1511.740 ;
        RECT 0.090 1489.340 2993.670 1510.580 ;
        RECT 4.300 1488.180 2993.670 1489.340 ;
        RECT 0.090 1466.940 2993.670 1488.180 ;
        RECT 4.300 1465.780 2993.670 1466.940 ;
        RECT 0.090 1444.540 2993.670 1465.780 ;
        RECT 4.300 1443.380 2993.670 1444.540 ;
        RECT 0.090 1422.140 2993.670 1443.380 ;
        RECT 4.300 1420.980 2993.670 1422.140 ;
        RECT 0.090 1399.740 2993.670 1420.980 ;
        RECT 4.300 1398.580 2993.670 1399.740 ;
        RECT 0.090 1377.340 2993.670 1398.580 ;
        RECT 4.300 1376.180 2993.670 1377.340 ;
        RECT 0.090 1354.940 2993.670 1376.180 ;
        RECT 4.300 1353.780 2993.670 1354.940 ;
        RECT 0.090 1332.540 2993.670 1353.780 ;
        RECT 4.300 1331.380 2993.670 1332.540 ;
        RECT 0.090 1310.140 2993.670 1331.380 ;
        RECT 4.300 1308.980 2993.670 1310.140 ;
        RECT 0.090 1287.740 2993.670 1308.980 ;
        RECT 4.300 1286.580 2993.670 1287.740 ;
        RECT 0.090 1265.340 2993.670 1286.580 ;
        RECT 4.300 1264.180 2993.670 1265.340 ;
        RECT 0.090 1242.940 2993.670 1264.180 ;
        RECT 4.300 1241.780 2993.670 1242.940 ;
        RECT 0.090 1220.540 2993.670 1241.780 ;
        RECT 4.300 1219.380 2993.670 1220.540 ;
        RECT 0.090 1198.140 2993.670 1219.380 ;
        RECT 4.300 1196.980 2993.670 1198.140 ;
        RECT 0.090 1175.740 2993.670 1196.980 ;
        RECT 4.300 1174.580 2993.670 1175.740 ;
        RECT 0.090 1153.340 2993.670 1174.580 ;
        RECT 4.300 1152.180 2993.670 1153.340 ;
        RECT 0.090 1130.940 2993.670 1152.180 ;
        RECT 4.300 1129.780 2993.670 1130.940 ;
        RECT 0.090 1108.540 2993.670 1129.780 ;
        RECT 4.300 1107.380 2993.670 1108.540 ;
        RECT 0.090 1086.140 2993.670 1107.380 ;
        RECT 4.300 1084.980 2993.670 1086.140 ;
        RECT 0.090 1063.740 2993.670 1084.980 ;
        RECT 4.300 1062.580 2993.670 1063.740 ;
        RECT 0.090 1041.340 2993.670 1062.580 ;
        RECT 4.300 1040.180 2993.670 1041.340 ;
        RECT 0.090 1018.940 2993.670 1040.180 ;
        RECT 4.300 1017.780 2993.670 1018.940 ;
        RECT 0.090 996.540 2993.670 1017.780 ;
        RECT 4.300 995.380 2993.670 996.540 ;
        RECT 0.090 974.140 2993.670 995.380 ;
        RECT 4.300 972.980 2993.670 974.140 ;
        RECT 0.090 951.740 2993.670 972.980 ;
        RECT 4.300 950.580 2993.670 951.740 ;
        RECT 0.090 929.340 2993.670 950.580 ;
        RECT 4.300 928.180 2993.670 929.340 ;
        RECT 0.090 906.940 2993.670 928.180 ;
        RECT 4.300 905.780 2993.670 906.940 ;
        RECT 0.090 884.540 2993.670 905.780 ;
        RECT 4.300 883.380 2993.670 884.540 ;
        RECT 0.090 862.140 2993.670 883.380 ;
        RECT 4.300 860.980 2993.670 862.140 ;
        RECT 0.090 839.740 2993.670 860.980 ;
        RECT 4.300 838.580 2993.670 839.740 ;
        RECT 0.090 817.340 2993.670 838.580 ;
        RECT 4.300 816.180 2993.670 817.340 ;
        RECT 0.090 794.940 2993.670 816.180 ;
        RECT 4.300 793.780 2993.670 794.940 ;
        RECT 0.090 772.540 2993.670 793.780 ;
        RECT 4.300 771.380 2993.670 772.540 ;
        RECT 0.090 750.140 2993.670 771.380 ;
        RECT 4.300 748.980 2993.670 750.140 ;
        RECT 0.090 727.740 2993.670 748.980 ;
        RECT 4.300 726.580 2993.670 727.740 ;
        RECT 0.090 705.340 2993.670 726.580 ;
        RECT 4.300 704.180 2993.670 705.340 ;
        RECT 0.090 682.940 2993.670 704.180 ;
        RECT 4.300 681.780 2993.670 682.940 ;
        RECT 0.090 660.540 2993.670 681.780 ;
        RECT 4.300 659.380 2993.670 660.540 ;
        RECT 0.090 638.140 2993.670 659.380 ;
        RECT 4.300 636.980 2993.670 638.140 ;
        RECT 0.090 615.740 2993.670 636.980 ;
        RECT 4.300 614.580 2993.670 615.740 ;
        RECT 0.090 593.340 2993.670 614.580 ;
        RECT 4.300 592.180 2993.670 593.340 ;
        RECT 0.090 570.940 2993.670 592.180 ;
        RECT 4.300 569.780 2993.670 570.940 ;
        RECT 0.090 548.540 2993.670 569.780 ;
        RECT 4.300 547.380 2993.670 548.540 ;
        RECT 0.090 526.140 2993.670 547.380 ;
        RECT 4.300 524.980 2993.670 526.140 ;
        RECT 0.090 503.740 2993.670 524.980 ;
        RECT 4.300 502.580 2993.670 503.740 ;
        RECT 0.090 481.340 2993.670 502.580 ;
        RECT 4.300 480.180 2993.670 481.340 ;
        RECT 0.090 458.940 2993.670 480.180 ;
        RECT 4.300 457.780 2993.670 458.940 ;
        RECT 0.090 436.540 2993.670 457.780 ;
        RECT 4.300 435.380 2993.670 436.540 ;
        RECT 0.090 414.140 2993.670 435.380 ;
        RECT 4.300 412.980 2993.670 414.140 ;
        RECT 0.090 391.740 2993.670 412.980 ;
        RECT 4.300 390.580 2993.670 391.740 ;
        RECT 0.090 369.340 2993.670 390.580 ;
        RECT 4.300 368.180 2993.670 369.340 ;
        RECT 0.090 346.940 2993.670 368.180 ;
        RECT 4.300 345.780 2993.670 346.940 ;
        RECT 0.090 324.540 2993.670 345.780 ;
        RECT 4.300 323.380 2993.670 324.540 ;
        RECT 0.090 302.140 2993.670 323.380 ;
        RECT 4.300 300.980 2993.670 302.140 ;
        RECT 0.090 279.740 2993.670 300.980 ;
        RECT 4.300 278.580 2993.670 279.740 ;
        RECT 0.090 257.340 2993.670 278.580 ;
        RECT 4.300 256.180 2993.670 257.340 ;
        RECT 0.090 234.940 2993.670 256.180 ;
        RECT 4.300 233.780 2993.670 234.940 ;
        RECT 0.090 212.540 2993.670 233.780 ;
        RECT 4.300 211.380 2993.670 212.540 ;
        RECT 0.090 190.140 2993.670 211.380 ;
        RECT 4.300 188.980 2993.670 190.140 ;
        RECT 0.090 167.740 2993.670 188.980 ;
        RECT 4.300 166.580 2993.670 167.740 ;
        RECT 0.090 145.340 2993.670 166.580 ;
        RECT 4.300 144.180 2993.670 145.340 ;
        RECT 0.090 122.940 2993.670 144.180 ;
        RECT 4.300 121.780 2993.670 122.940 ;
        RECT 0.090 100.540 2993.670 121.780 ;
        RECT 4.300 99.380 2993.670 100.540 ;
        RECT 0.090 78.140 2993.670 99.380 ;
        RECT 4.300 76.980 2993.670 78.140 ;
        RECT 0.090 55.740 2993.670 76.980 ;
        RECT 4.300 54.580 2993.670 55.740 ;
        RECT 0.090 0.140 2993.670 54.580 ;
      LAYER Metal4 ;
        RECT 7.980 2983.720 2989.700 2999.830 ;
        RECT 7.980 15.080 21.940 2983.720 ;
        RECT 24.140 15.080 98.740 2983.720 ;
        RECT 100.940 15.080 175.540 2983.720 ;
        RECT 177.740 15.080 252.340 2983.720 ;
        RECT 254.540 15.080 329.140 2983.720 ;
        RECT 331.340 15.080 405.940 2983.720 ;
        RECT 408.140 15.080 482.740 2983.720 ;
        RECT 484.940 15.080 559.540 2983.720 ;
        RECT 561.740 15.080 636.340 2983.720 ;
        RECT 638.540 15.080 713.140 2983.720 ;
        RECT 715.340 15.080 789.940 2983.720 ;
        RECT 792.140 15.080 866.740 2983.720 ;
        RECT 868.940 15.080 943.540 2983.720 ;
        RECT 945.740 15.080 1020.340 2983.720 ;
        RECT 1022.540 15.080 1097.140 2983.720 ;
        RECT 1099.340 15.080 1173.940 2983.720 ;
        RECT 1176.140 15.080 1250.740 2983.720 ;
        RECT 1252.940 15.080 1327.540 2983.720 ;
        RECT 1329.740 15.080 1404.340 2983.720 ;
        RECT 1406.540 15.080 1481.140 2983.720 ;
        RECT 1483.340 15.080 1557.940 2983.720 ;
        RECT 1560.140 15.080 1634.740 2983.720 ;
        RECT 1636.940 15.080 1711.540 2983.720 ;
        RECT 1713.740 15.080 1788.340 2983.720 ;
        RECT 1790.540 15.080 1865.140 2983.720 ;
        RECT 1867.340 15.080 1941.940 2983.720 ;
        RECT 1944.140 15.080 2018.740 2983.720 ;
        RECT 2020.940 15.080 2095.540 2983.720 ;
        RECT 2097.740 15.080 2172.340 2983.720 ;
        RECT 2174.540 15.080 2249.140 2983.720 ;
        RECT 2251.340 15.080 2325.940 2983.720 ;
        RECT 2328.140 15.080 2402.740 2983.720 ;
        RECT 2404.940 15.080 2479.540 2983.720 ;
        RECT 2481.740 15.080 2556.340 2983.720 ;
        RECT 2558.540 15.080 2633.140 2983.720 ;
        RECT 2635.340 15.080 2709.940 2983.720 ;
        RECT 2712.140 15.080 2786.740 2983.720 ;
        RECT 2788.940 15.080 2863.540 2983.720 ;
        RECT 2865.740 15.080 2940.340 2983.720 ;
        RECT 2942.540 15.080 2989.700 2983.720 ;
        RECT 7.980 0.090 2989.700 15.080 ;
  END
END SoC
END LIBRARY

