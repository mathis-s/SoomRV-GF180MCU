magic
tech gf180mcuD
magscale 1 5
timestamp 1701464064
<< obsm1 >>
rect 500 500 43686 48988
<< metal2 >>
rect 1872 49188 1928 49588
rect 2222 49188 2278 49588
rect 2672 49188 2728 49588
rect 6722 49188 6778 49588
rect 7072 49188 7128 49588
rect 7272 49188 7328 49588
rect 7497 49188 7553 49588
rect 7722 49188 7778 49588
rect 8022 49188 8078 49588
rect 12122 49188 12178 49588
rect 12522 49188 12578 49588
rect 12872 49188 12928 49588
rect 15472 49188 15528 49588
rect 15972 49188 16028 49588
rect 16372 49188 16428 49588
rect 16672 49188 16728 49588
rect 18422 49188 18478 49588
rect 23284 49188 23340 49588
rect 26472 49188 26528 49588
rect 27322 49188 27378 49588
rect 27440 49188 27496 49588
rect 27664 49188 27720 49588
rect 28172 49188 28228 49588
rect 29622 49188 29678 49588
rect 31672 49188 31728 49588
rect 31872 49188 31928 49588
rect 32472 49188 32528 49588
rect 36522 49188 36578 49588
rect 36872 49188 36928 49588
rect 37072 49188 37128 49588
rect 37272 49188 37328 49588
rect 37472 49188 37528 49588
rect 37822 49188 37878 49588
rect 41922 49188 41978 49588
rect 42322 49188 42378 49588
rect 42672 49188 42728 49588
<< obsm2 >>
rect 500 49158 1842 49252
rect 1958 49158 2192 49252
rect 2308 49158 2642 49252
rect 2758 49158 6692 49252
rect 6808 49158 7042 49252
rect 7158 49158 7242 49252
rect 7358 49158 7467 49252
rect 7583 49158 7692 49252
rect 7808 49158 7992 49252
rect 8108 49158 12092 49252
rect 12208 49158 12492 49252
rect 12608 49158 12842 49252
rect 12958 49158 15442 49252
rect 15558 49158 15942 49252
rect 16058 49158 16342 49252
rect 16458 49158 16642 49252
rect 16758 49158 18392 49252
rect 18508 49158 23254 49252
rect 23370 49158 26442 49252
rect 26558 49158 27292 49252
rect 27408 49158 27410 49252
rect 27526 49158 27634 49252
rect 27750 49158 28142 49252
rect 28258 49158 29592 49252
rect 29708 49158 31642 49252
rect 31758 49158 31842 49252
rect 31958 49158 32442 49252
rect 32558 49158 36492 49252
rect 36608 49158 36842 49252
rect 36958 49158 37042 49252
rect 37158 49158 37242 49252
rect 37358 49158 37442 49252
rect 37558 49158 37792 49252
rect 37908 49158 41892 49252
rect 42008 49158 42292 49252
rect 42408 49158 42642 49252
rect 42758 49158 43686 49252
rect 500 500 43686 49158
<< obsm3 >>
rect 500 500 43686 49154
<< metal4 >>
rect 522 1568 822 47824
rect 922 1568 1222 47824
rect 42863 1568 43163 47824
rect 43263 1568 43563 47824
<< labels >>
rlabel metal2 s 26472 49188 26528 49588 6 A[0]
port 1 nsew signal input
rlabel metal2 s 27322 49188 27378 49588 6 A[1]
port 2 nsew signal input
rlabel metal2 s 28172 49188 28228 49588 6 A[2]
port 3 nsew signal input
rlabel metal2 s 15472 49188 15528 49588 6 A[3]
port 4 nsew signal input
rlabel metal2 s 15972 49188 16028 49588 6 A[4]
port 5 nsew signal input
rlabel metal2 s 16372 49188 16428 49588 6 A[5]
port 6 nsew signal input
rlabel metal2 s 16672 49188 16728 49588 6 A[6]
port 7 nsew signal input
rlabel metal2 s 27440 49188 27496 49588 6 A[7]
port 8 nsew signal input
rlabel metal2 s 27664 49188 27720 49588 6 A[8]
port 9 nsew signal input
rlabel metal2 s 18422 49188 18478 49588 6 CEN
port 10 nsew signal input
rlabel metal2 s 29622 49188 29678 49588 6 CLK
port 11 nsew signal input
rlabel metal2 s 42672 49188 42728 49588 6 D[0]
port 12 nsew signal input
rlabel metal2 s 37472 49188 37528 49588 6 D[1]
port 13 nsew signal input
rlabel metal2 s 36872 49188 36928 49588 6 D[2]
port 14 nsew signal input
rlabel metal2 s 31672 49188 31728 49588 6 D[3]
port 15 nsew signal input
rlabel metal2 s 12872 49188 12928 49588 6 D[4]
port 16 nsew signal input
rlabel metal2 s 7722 49188 7778 49588 6 D[5]
port 17 nsew signal input
rlabel metal2 s 7072 49188 7128 49588 6 D[6]
port 18 nsew signal input
rlabel metal2 s 1872 49188 1928 49588 6 D[7]
port 19 nsew signal input
rlabel metal2 s 23284 49188 23340 49588 6 GWEN
port 20 nsew signal input
rlabel metal2 s 41922 49188 41978 49588 6 Q[0]
port 21 nsew signal output
rlabel metal2 s 37822 49188 37878 49588 6 Q[1]
port 22 nsew signal output
rlabel metal2 s 36522 49188 36578 49588 6 Q[2]
port 23 nsew signal output
rlabel metal2 s 32472 49188 32528 49588 6 Q[3]
port 24 nsew signal output
rlabel metal2 s 12122 49188 12178 49588 6 Q[4]
port 25 nsew signal output
rlabel metal2 s 8022 49188 8078 49588 6 Q[5]
port 26 nsew signal output
rlabel metal2 s 6722 49188 6778 49588 6 Q[6]
port 27 nsew signal output
rlabel metal2 s 2672 49188 2728 49588 6 Q[7]
port 28 nsew signal output
rlabel metal4 s 522 1568 822 47824 6 VDD
port 29 nsew power bidirectional
rlabel metal4 s 42863 1568 43163 47824 6 VDD
port 29 nsew power bidirectional
rlabel metal4 s 922 1568 1222 47824 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 43263 1568 43563 47824 6 VSS
port 30 nsew ground bidirectional
rlabel metal2 s 42322 49188 42378 49588 6 WEN[0]
port 31 nsew signal input
rlabel metal2 s 37272 49188 37328 49588 6 WEN[1]
port 32 nsew signal input
rlabel metal2 s 37072 49188 37128 49588 6 WEN[2]
port 33 nsew signal input
rlabel metal2 s 31872 49188 31928 49588 6 WEN[3]
port 34 nsew signal input
rlabel metal2 s 12522 49188 12578 49588 6 WEN[4]
port 35 nsew signal input
rlabel metal2 s 7497 49188 7553 49588 6 WEN[5]
port 36 nsew signal input
rlabel metal2 s 7272 49188 7328 49588 6 WEN[6]
port 37 nsew signal input
rlabel metal2 s 2222 49188 2278 49588 6 WEN[7]
port 38 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 44486 49588
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3136006
string GDS_FILE /home/m/Builds/caravel_user_project/openlane/gf180_ram_512x8_wrapper/runs/23_12_01_21_54/results/signoff/gf180_ram_512x8_wrapper.magic.gds
string GDS_START 2941552
<< end >>

